��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$��4�o;�����~>fF��i7����l`Û�%�l{t�r	�@Em�,�B=���Z�Vi�?�v��P�U�=�
��ۅf����u��ɡJמ��+"9e)xpƱ�7���r�CƖĽ-�=fK��ٞ�yq|J���\���t��(�B�^�=�S���Ȝ��܊6'{�߯AI.a��`=uzmu��g\'x𺼕�͢�*�g[+�CwT'r���ӱ��*��[��B�g�d��׌w���G��2�ޚ���l��k�۸�m�i(b[�{�㇌�]�i�5'�`;Etg
<������H�W޵α�𧝅=��q·�{���TgU��tU��Y�ʶ�Z��P�[�8�����,���3[	���@?���8�?���A�ڻ���xY&�a�Yz�t���8S�
�t��'�bh�V��˅��:Cf���Ì�{��޳�`u�p�Ө��0*����� �ʿ3����{V�dq�M��gP03�[�noܫ���wP��HO�rd�v��(���?���yk=��\S����:�\���$�t߶��+ދYk��},d���`9 n�>�`��}}�"%�zR��B[�ήN� ��ǜ׊��&*]'����tS-͐!(�������_�Qj���X����N�v���B㷙��ٍ��\T��1�ޢ�͛��Tߚ��n:�ň޸'&Z��~3#$o��Q-�%V��172�==�u-[UA���'89�g֒f�IY��"���ϙ����W�8��x���+�yO��s�Qٴһ)>`u-b��C�I%O.�|PB��[�S*!;i�U�Q��m��E�0���|S�{J�vX������`Y�N��2r�m�JO��[}��T!B�S�� ���|^����n�ᐧ�������"tC�]���;�'hoW	�4�G��-��L�GD�5���Gg��n�|#B�2
�ܸ�b���%i*dH|�@��֯""+���S&�'�{3V�8y��r+��O.S����E�$��0�������щ�.��\�4�?����ޖ��ŵ��-����G��!�<���'W����}�	�73�")9�@�/(q�~� !�?�O`PA{Ӆ������'�b��[S�����|n8	n�VGB,��-�[�>;[tm�a�&�E<V�ɎӜ�������.��]�Zut���e������Ԋ�1��:��s�X��jt&��2�ĭ𧦰G٭0Y�XZ^.���)��q�t=7|	6��$�"����'�>�}�e�~���2r~£^z;��J�.��BuӋD�&�u��`���	3P���;��o:V�i����i%��H�h��)6��8(ξ�L��u��q7	�}WɯP���������$yL�ڠ��p�k����F�;�G�8�,� ��`�Je��O�B_�=����/��L�>t�)9���9ތ ��ey� ����-fr��Q"^ b�"כ�m���~��.;O@H�~�;sN�x:�a����� j�y�_��pZ<)W�N��_���9z���vÄ�����䫈�cȸ�o>x��1��$&(:!���v`��w����BCr������}9�\��9`M��Ǽ�"��r�����;�\q��Q_���ɖ�ώ� �ϩ�:2s���C��- ^� B���S�W�= >�}�}(9�s.)U�h���BE=��S"o�D�wF��	Բ|���i�ӏ���¢6�����7z�d��`�I+0�/E��P���6��-휒�N�)��Mߐl����#Cؖݤ\��'^+NЗ>Ô�(�ԃU#���Ϣ��~�,��r���B92���wQr·_`�+Ux���S�o2l�*��Q���>��t�ɛ��e��A�B<$��~�.XZ
p�<��㸇!��P��Sf֭�7�X��IN���:]���"�O��A�z�*���R���x����2�2�)�H��mfg:�Iv`X�in("��v|�w?2v�y��q����]�C�k�_2c�&��{�T�p �j�n�?b-×�>�|)u��-�k$��eW��0�z f�aU�Jg�,'��z��ͼb�sX��FK��� _䧙�eQ�2�jf>�K�!�C��{���n~2�I(���A�~A��<�]���e~Q��vR쓎�j3�r��]O�"��v����VJb!ǅ�fF�Ҍ�k�
T��1)o(��q$y����W����i�������Zv���B���Z�)�s��yo&��C�N�^�<U��� �IIP�
d��\�o�M�[r��>V�9�4�+�Q�}�h^��´	���׵���&�3��4���#�^�Y�OU�h�;������V����9F�c�`\�[j�Z�./7�>0�9����0�T��yB��EU��������p�	R	T+ �f����꯯R��v@#^�h������<����i��=)2�13 ef�I�\;	R�[�6��:���%�;/�`;ϛ�OR��������zY�g��x1��|��A�m�`�Cp�lŔ�N1z��A]��i@ڄ���f�ʔ�ė��oss/�|_A�;It� �(=FF!���H%Ȃ �V�y^�J�!�W�����&C6��㐙N_�j�)�;�V$?I����W&�Q���D�,O�K>D����7��:Bo-��y+�>=M�'��;�H�?4Խ�<�j��ucW�.��9;���H��vw9��Fev{�)����`G����R�k���p��X�S������W�8{q�\����D~m�'�0�}�9�L�%�
��p���<�x��{��C 9#�!�1�o�-��+҃�=����e��f ���UŻ[�̺z��L"��	n�@��"��:�j��X��1�-x1�v����\�u;�'�}JT|�=Էn&b�֚_�&�+)�t#��H��� ��&�9m$6�K����r8ak{�����?��S�:��f^�Ml���1+�Ũ ��7��A&��D���V��E����/͉�8�)]�ZW9�|m >�
�/�U�Ѓ��S�,\�ĕP�x����D�  7Ř[6���W�T�[���E��,��s�w	}�2�`1��n�� ��D��ME��>�${G���\���5xj� (p+�iTV���R|?co�_�?o��a+�q��I��E������I�Eθ$#��e0����,����|���y�%��II���`���t�;�A��&B��J2՜���|�^E�F�FW������=Ǹ�
�%
6��c�n9ֻ�#O,ѯU�K�:����A�Q���+و%~�/s�_�U��I���a@���O��>�����ȼ�R'������0�FUQa�8�D5FcO}�j���1:���������2[��c�;�J�8���^Ƽ�si��\���[M��� j�	��k�2ş��J��IK�~o��q�Ol��BQ��2�CZ�)�d_�f�����b����N?�:C�9��/[�-�?�;fn����G�����-�W,\f��V�OؐO__��/u��2
���v�4^��)j^v�IU\��}3��&�俁��&�4Hi��.M��,�5Y�����1c�>F�B���{�Z��&Ύ�:]�,������&�q��6xa%Y�w���Q�60�xC>T��g���<v����&�����ohP��.���a��Zb0[�yh��ˣW����M�䶤8nW���٠�X�m؆TO�OH�R�=����p%�/�>l&�J�r�D�\�"���Ylt�H]�<��'��\�xq}P\�J�e$��Q��۳	B�|�e�@-!��3˷v��6�.1�L"��(��ው��q���po�cs��q���)/�Kzs]=����ǗMp��QR��'a�M����i�����-���p�q25lq�t|�Y������1��c�	na�=�7��fE�$��wܨ���忹ǤD3��s�A~yu�|��3�{�V,k�UvVO�i;e�0H��W�ͫ�{܀ی�8�y�"')-vU�s
>H�Z�${���Sz�
��<�J��n�k�����$����"��%��nb�']��cg��^�uڦ��)vɶ�^��6�U�3���Gw(��t~��p�����N�P�7�'�L���k��`�Քаc�\^�dW�p�Yd��?e C~�;�b���,�:�^$HYc��{:�rt�����m������6
��q�ͽƸ�ȉ��I���8Z��J`t�!VB)&��m��@��uL�Ҟ�n{	s��$ԕ��§\�p���R,�O�S2+r�{�Չ�䨳�4�� ;ӵV	����E�R��?���.bOd�ljr �{��vvf�H(y�ٮ%�Oи>�"�d+����A�u����_�o�V@�|�5j�*���FZ��V$�I�I�w咲G4������gk���G�����G��#�V�X�ߋw�q hp�6S8�H�ܰ|-���<X�Gz�%��opv%:�f}l_�9'T9Sյe�(C՛�n��޿�oQ�g�#�����N��є0eG돽n���7Etc۰%n%�C���D�pȥ�C�f�� 'nm>>}a��%n
W��f��r_eh�3�bG�:[D�P���Fn��}$�v�o~9[�p�f{�[���5Ey4�&,�"���!2-[8������� p
N^�G�}����W]$zv�cҪ)pR&?���Y�Yc R�a��`jc��k�<�8���!�̍�֢�<�D\�ݦ}�B��f���F����zX@(�<6pҕ�j��shF��+̚HtKV!���LSv�E�^�&1U��e+*�c�s�,g\��[͸�\�[�S�ҏ�ɽf��RŃ�:�g����<�4]zd�[E?B�c09�{��il�*I]�*�2�yԷ6R|��4M.-�]���@m{�ي-�N�Nƻ,��ƦxE��񤎘����iZ|,c���?o��Y�Le�Vz�0-_����%�֪T�R��4xV�C_��0ÍHs��n�0~��N�����n��cФr�3G�~M֮��\�j���S��cF� BK�q�C��=��S��-W��Sy~p���:� ��
c�-Z����×�jSz��C^�[
L;kN�m܁�x,1d	���d�����0]�l�m�L|y/&�z6ѧ�����b"b}����C}8R,=���)/'����S^#ҳ���Jn���$��q��hvQ���1�:L^����N�4�T�!�,�����8ӆ C��DS��3�d���\1�l��
s��{��:9f0�)��.���;sl�a�1D]�j�4R�Sg�Z���8I6�� 7�+��_���Y�>Q��p�}񬛅�9�G?��,ŷ�-a\���I��L]�F�1�>8:��\�9��n��|긲o��o����#�Q!�Pǋҳ$��E�\~��_'>0��X�{G"���I]1���2��1zE�3a�W�SZ8pDKC�*���qS4�i�){���g����U�Z�f'�X;a�9�Iƞ��wMT����N:<�6�Y�fz�j!,����E'��QmR�\^�_�"�8�4���)#ʧ�3�u!Wi�۔�~R&�	�$�n��$����fZ�c��9�^�pi�x�T�$zzO�{L���r���l�䃝v�r��D�
��P��U>,����b��f�<@O42��s��eS��"A�����R7�C�B���5E%�{�����T4��C����z)ɋ�¹�!H�1�J����lar�R����;��4<�i�<�%c�Aœ���\�c�7Vk
?� W(��ib�-�y��=Ծ>P,�L]�-�6'P ��P�Rb1L����=��!���>=_�;�r�wRH�Q�h�p>v�����+������I���~���s��`�ڄtU-�{8�+�ȏ�3_�_ų�w�Z�_n��[O�C�H_���?���x�川��c9.��O����``�=��ǝ�(3��Eɻ��>Ķ͒H2,����s%7���w([��Zt���ຄm�l�˂�ea��+�^)/��Q6�#g�t��}�YN֬� ���:����4��*rخ<&��'���LSe>��$�yPMi~��6�0���Zʞ�N�P:���y	t�f;�um�W��������%-���Ȥ	�T]�k�O|�C�='�l����ۗ練|��b�6$T���sz�[�AK=6Ŕw�śv��F�6��&'Ϣ&L0uc_F`�Cº~��Ss����0t�m�C�T�T/�+Ȫ�)�Ar�+�B�e�T��U���O���բ�T����aa�7@Y�ZE����k9<U$?ZP0.�T�N1��	�~�z��h։y���e���u�=-��XO��w׽'o��@��4K�W��N��zN�mk���*������@��J�����ߍ����V�����a���t�h{��-�
g�\��^�Pp���3��싂UU��e��!I�-1۽��ե8�MT���Ԩ"����]Jnon���#�W �������W.'E��g�
�e'$g��ߖh_�a̕(�~U���T!��OV�p������,�����9$�� ��
a	����^Q�֔�b�Ӌ9���nk3�~+��TܕE��|D�*���8?�FD�k�nٟ�&0٩i5�1�R[� ��	8J0�|���w���+&��f@8�]6��1B�R���_� ��u�p�1�k��ϕp����}5�d���z����=�6$sd���������'�w�NG�����F��'����(/ņrv�{�D>��#��pw�ذj�K�����{~�@�z,5wጸ5X���������S����ޅH(MJlO�S���k̟)�؉��!�J{���d�5/
n��~�^i�>$�H�u��?)YR���6�w�������t�l��Gaz�}�ⲆIǠM̾Vz��@(���gD�Xg�gʳ���Y:$�	���x�YP����HH�ۗ��/(A//��i�i��D�I�"?1���3�S8�+���%F�K�?�%���~��5��/�u����[�9�������Y*�y�]�RMD�'�aTMU\#�=k:D�k߬�uF��B)�3L[��@�xPk�����s"�+u�$*��/�4߿��Y�!�~����^$��NM��~�77�՘qjc=�z�|����^1�.\���xD���1���ug�Rza���:�*�S���
��?g4ަ�S%�6�U�����k]�0��K�YF�j��`�oaž�+>v����gH������{ett�p�,��G��k�bs���њ�l����lj��C�����<Y?"t���=�=aq�7�?��[d��%*��5(�uj-�Xe���D�6�wW ل/г*��}�0��<?3!��A���B_�U{�� P;ܔn:����kJ�לr�ڢ��ӥ���4���qZ�Չz���՜z��`WS�SU���� 8&W $v����ri�c4˹D0������	��1�*�-T׶\����(�u|i]�P�&���f�6���4£n���n��L]k*��\�d��%y�E��ب��/hT吰S��V0���������'f�_ê���`��tm��;kvy��&�����}�׸��OzA�\��C]\Z�)+?�6c�"����Z�H�۞1L����4A[�]V�w-/֚C�P���¿�ae�C;�a����� ���$�r;��o �'[����V6	�Cb9��PM�`�Kc�{lF�܃I>�Is���$ܱQO ��-nH�a��l8!�[	�0L��)��;�Yp�E��Իb��]�Vܶ�𭹲����$��*�L�:(YbC)�v���YQ*��������-ʮ1!`��qHai�p^x�z�Q�Qp~�0R���?�ۛ����^wH����ݝ�Gd*�q�����T?������G�.F��F�+�ނ�5��'˻�����!I*��&�^)Yv�]�h���X.d��� �M�f�� ��IвМ�K�55���������UG��0N�� �؈&
��#����bE�.2ݱ�抱�ueC�	��k��>��e��\\:��9VN};J����Q  ��O�k�)�o�U�\l#��G**���l\����������rN�u.�97�⿜�EN�V �~�|�Nv�j�aVq2÷��p��1�T�KlO���@[Hw��lY!�H�<V!<?-Tn����\<�s�@<�9D���G�?��r�M�
+IT�����n'�z�5
�o�Ʀ1��������s{�0S/ft$����@OtXԳ����]�
����J89�0OzR\P��S�g�v����a�nCrߖI_��h�)J�Y�|��,\��[�}��h4}�%zNE��k�R�����g���>7���I+������Uʜ]yLK�%X6<��f��Gd�!�I�M%��\��Po3�I�y���B����jИ-xJΨ��~E�%~lw�؈���56�T��R]�f	���t�k�`d��F���lkШ �=\Z�EC[i��G	ᇢ�E��{Z���������O<�%T����p��t�2yls�,�Z��6U���͡�2��(6Wi�u���z}`���7�� �:����O[%
&�gz�'#}�u�(��\�RU�ˢ���]��m,1#�r�=Pׯ�+x�r��y��޽bNl��),I:4L������l7c��q�Um'=�m���q��x�ǲ����+��#/!� }3!�\u��9���B����0d	�8��`>�7�3/Ml�](���������E�S���=drOР�)aiQ�t��S���*ط�"��/��{O�5F�}[�R�G����;72��@֊H/�
~��;�����8��r(
󟒻�0��l��|M,=Ք=���H����>�fw3�=#54�l�ZF��T	�G�$'�J����X�/,����Q�5��S��=׮lKC���c�J[K�]n����hO6k��j��_Ǹ�#��pe����J|��UU?L��`s&��3��ؼhT��e�����$,(L

~���w�N���M0K{�c*��0����1��
-�Y嶂26�;�c`e�:j����V�-��Nc�iL!���a���B)�pǉ$4��`qT�ٲ�e�<��eQ�)��F�� �+��o�J|�C�/�Ԋ�d4@���?&�%�.�|a����!uo���m�tJi��f(��'��8h�,-O���d;��@ݙ��]��:,��nIt��ʀP�x���o$�c���.KU4�8�p<����Ɇ�k�z`��Nͨs�:�*�x�t�����p�����j�����K�}�H1v���<7��V`�4�u��X���?4U����8�
n�Ei�*��.�Y<���26#Ƨ(���)<-K��x�sJ'&CSF�p����@�t��-�{����%������@L�^�g3�y�$�	��An�׮�r�Pk�Q~Ǻ��~8�<�rl�#��9��X�@��[�; �uɀ����'w���D���j��×��]L��v���ꄛ<�p��U5(�c1�q�y�z����U˒���
���;�G,t<�7�_��c��`RQခ���(n�������@U5�J�5O~�j � �ԡG���}�N�k�vY�20|*�`����"V��H7M��m)��a��0��f=焞e�����`zǔ��!.��@D��3�xR���&T<6��/�>�cM�M�aJ$�>v4�r��Q�(�eX���K6]Ub�*O�}{y�ɍCW��!bb��+��Kv�����7��#��^]�&�z',Ըn7�����%�gR�B��!�v
��.���7�A�Ҷ��D�t?�p��Te�\���e�i�ˆ7#}C��_+�'����8��i�q���7�5\�[��O��v>�V[.�m��e@�R����^2��(M3'8V'�q�(��?1t��P(� Ka.+)������,jo����PSL��wBZղg���1S�ᕒ��?�([��,�hl����*�-�w��/@�5UPr�pl\2ueL���B��Tw���Qx���wJ�9�!I�9��!h�N�.u,�Ǳ�"����m!����J�pV���䁓��;�k%@�ZD�$�F�!�7,%��Ғ������z�����]m��%6��#5�4���y������Ǒ�Xc�����<٤�8�8;���O� �hmR�O�cW2Y��q�}#��mN�;���1�J%q��N֥1�����g��M��,T̞�W�mHi�@:�&�����~ZG�~���������j��'��Ff�e�ٵ!Őa�������u�V��Ib��NK:��sN�o�����l ���Q�Ay@�X�>;�+s)5�a�JЗ
��[�?4_���Y�'�R憁�>�ʉ�yrD��"��ɟA�kLӉ��BׁD�"����n��\��^�zik����<d$�~u����2��KCi�=���Z{���w1>5�JS�WТ��wZ���1�Ykc~�.�����^�CGӇ��M+B6\��/��	RC������	�Q�w�A��`�����J��o	%�؛=�����鑬�m����7�5v���]�ڢ�lU���i���yGU��ǽ���.�� p��h�6E*�ܧ�6`�����-��c>�9��x��a��呼Cm> T]�ly�E�B@\�4=٭��36r�6���d�;<�))��鋯"@}�DZ�CI"b�#'���h"�L�� e�ɵ~&p<e��J�(��.�Sm}��[���?�Q�P6)�u��/-
yX�-6Rdi��~���i���.օ��	d��c֎�Cq6��AT��,Gep��.������"7�&���{?-:�O�*q��m~zq��]'��!�_�q3T)!����ⷔ�π0bIU�-���[�UT&Rlx�85w����N�b��bUF/0��-������q�$OW0u� �%�&� �Nl6c�D��Z�������	��	�1��k̆�{=�yl��?������ظG�א��o'�>��q�G�o��H+�����9��3(A��p�����jT=EP�˼BO�{�TQ�~yU��*ɏ�õse*�yy
���-�g�z(�_�1J�O�&�.ϺB����
*��z�H��b��-�/�$�V�5�z��ժWD囧*�݂���$�W��H~�Vte�*��l�|�����[�xG��z�'�Ig�\�X�Ka^�1���/!ֶ����c�&�X����|Z�,�F�/dy����R��F��~c�D��L��'�xݗSN�_|,ʋ��Za VOe� �\�v� a�L� ���0�l�ˍ�OE;����m X�L�����C1}��	���[�o���X�%l
;��UUэN�fS��e�L�B���܉���ǣ�k� 2ce�`�����-�����e��,Â �μk�|�P:�*u������Pt�8Τ`�ڴo�(���dG��.��(y�WؚK3�����o��'��wvNY�z`f��>iv�e%f�FW�c2`�(hH�}+jm���kr{ E�@�o'	
Ǖ-T�4lQ�XV6���'��f��L�U	$����EQ5�A�Xe;�44��=q[���l�5r�G�\+[��O�l_�����x��c:ӑ��z:����v�����p��2��V�^?3x��y��5��ʍz<d'-u8U�uݟ>Ig���:e��O^Nw}z��ڨ5]�j"�tbdɺE��R�Q|��a�r#E���qx���%�V��a<��-v'"�F��-�~���X��o�D�w�cM����ünl��!,��:Z��FJ��s��R��=�
8�H=?nK��Qz��ɮū��\AʰG0�%*�����<9�O=V����=T́1-�7��դ�?y��a�^�ԭT2��J�~�+�=��[)��T�g����T�#@FA�]��>�\̭��}\H��wҗ�o�,�����Q�#�,@�6�t�[����0��g�C�����L���WD�
8\`Y�g��p;S#j�/֝P͘ŴU���P˙I���A��O	>�.��� ���p"����M.(�A����d�^�Mɠ����1���n2�?�F�O��`�]�i���U����_��;��m��v�(��|���� ~~�]<�OKD�J�ob\�IF��h\�~r�Xʮ:��]WK�@�F��S�����\^_Q35CM!��p�媲1���p�]0}R��5���<O�ц%x�D�˾�ߜ{�A��8�����S�8�Y�>��嗷�QLS�u)�
���w�gFRYë��m�nZ%漢���b��\�6<Q��������W;����gE���r�n ��}6W2�O�  ��v�/�v���u1_�w;�t[�&�x��k��u<Gykߟ��a��e"G�^������H4�Gd�ʨ]���;5��Y�Rt��N�^���;��h���ZA�%�y7]��M��fuQ�I�^���6��iE���@�?z��k�ꚬ�c-�K��q�yXϦ��b�aŰ���*��o,j*��ls�BZ8�;�fդs�l�V�l��v|�YC��Ā�� A'�B�3� ����P��d͒)�Xȓ�hm�ͧK��o$D�VТ�a��8>��4��>�ds��/|?)u���|�,D�7��{c�vK9����)-�<�Ct⺅ se�5}�@�v����贊���bP���>�jI��[p�)�l��	$��dރ�w��Ҁ�-��dh�d�s��DW��Ń��D��
��oɇ���"��Ҁ���vr]ȶ5�l�	(����]���'fv�Lţ���=��34�f��[��"�rM�����N�+�(wY���ZC�r�2��fB���`U����ܚ����5X�T@�sn5 ��+���{�F�_�V���,��.J�Q�-H8�e���I-��&(EOl����Ƿ5��-�n�A7���⺡2s@$�ư�HA�N!009�TS�l�{��W�$����ٙ,>b��Z�Fx�"�sX�h�e(��G���ƒ[̏/�M����!�5�B��pĔ�&h�ƒ�O�q�K�jbfd?�7��x�M��Q�~�X_'F�{�Q��=��4y�Ǔ}X���1�.�Qz�N�Q\�^--�2��Z��������9���"��u�BZ\K��U#�bx�?���u��FhQ˺C���t^BfN!�U���Uv�w�?&(ׅ�$��>���:`QW�+�iW�a�t�.L�h��y��n�"5�SJ@3V�Z�P��^����M����]a}@^�=�6�g]9��C�av#�D xgaS,ݶ���),��G�z�[�+��|����B֋, ��l��'U_˼�1�m�����"��T�"!�M׻�����F��c~<�[g�h��_`�cF���9}�d��v�����H�c�a���s�biWd�!U�:����?�Ë�*�ۉ�~	Pp�b�9 ���F)�}����s��|(I/k5��_`7�'���u�& k;����aKŐ��?�	޽������J�5�x�Ƅ� �!^t� Q=������1$.����%�풻��iEZ�V�)��g�q$�|9uM:�Z;���h�+��W�+2^�*���8�;����n�OJ����	��U���j�aʀ<�޴�/F������h稛�~TP+��#1g�B�����;�K��S|%�b�D���`��@J2	� k���؞��S14Y�!!��z̊/KG���=nELJ���p��<q���v������Y"�ݱ�ӳ7��GmJq�A_��!��w�	�?1��D�
����fXE6�L
n���#<��x�ه	A�GpJ	��$�3]ngOw(	!R%I1����0箮�b�Z�*zո&�Q �}�s��/���~�4&����?<��5�އ_lW���z��L�@��|4�E/4߮�N.J���Z�u�;Ϥ�������{�d�L�b�$�fk����-R�9*��rl�r�4�%ԝRr�r�o���W`/+��eO���^�ۮG|+��g��S 
㱎F�FigЯW� ��I���H�����GPQ 5ߏ���4bRr���8��O�"8�v6������A%2W���l�W�OQ���܅�ш�i�xR[s��&�K�����a;6�_�!;��Wz�W�\�F��ɨ��QVq���ɍ��:yA��N�乑	�m�G���(���d)��]J��,���,��j{�r-y��Kd1����/-���b3�3&�9,�b�GdK��B6���o�Yo��Ql�b��9#4������#$��]Q��{�3
!mb9�(�H'��jt��?K�,�L�*�4���Q)&\�?��Ć�1��PJ%��[2f�(�]�`�iﶹ�̈~�d����4�Y�/�-VPܔ��.�a�]�[T��--�cEuf�S���l����ސ���6��=U�����@H���Q@	J�����zd�����-�V�ǈ-��vDU��.E�0癣ڲs�}[����mYE����.Kp5��{˼a��MO�Yр{�Gt;�n���@��x~Ëu�.��]�k��0n�2\�3dAJ�9��x�8!����L�f���J?bݷX@?�I���p��Tg�ف���:�����gӂ�م�˰��&Ƙ��t�����|S��7�=����RT39L�	�������Y(�*�F�d���K�`��@�q�0-x��MZpE�,��Rj�XĻ��U��(�%m>i�~���C�YG}�(~D$6u-����DL�/l��N+g_�u{�������-�7d0�T�S�c�\q.��56}�V[�c�~�,�v�JK�udQy���e�g����[��s�(�5���6�湟_{��預����@i+a�ds��P\&�1�N����+��I{d�dPK _X�uqy$�k����6_�*�$��NH��<��D��J���Wu�x�d���1�cTA�>��v��jZ�̟J&�_ ���{�r�C�������C"�(B˱�a��+�h �1J/v-q<�-�/ۄ��0���ժ�N5�/���%5�L�8VO��6
 kkCW�Wm�P3�4�WF�_�3c�E��Do����)��!�#3�"O��GU�>�U}.l��ʹ�3�w-x+k@��
}�f2�Ǽ��ǡRG�}r�M��	)��C�ѹv#˶s�����~A�a�����Ӱ�H��豜$vHXgL�iy(X����;cm�I�&�0��9X$�������k��'���<j6�s�!	w�N������J����K{O�M̈���]��;I�!��bnד,���ԑOn�#!	�B�qL�z����l@�����m���V����R�Y���)��W�G΍ϯ�������t N1�l������D��.u��T5
^��J��~])�P�J��s�m/�-���0 h��J����|�g��Fo��+���7��i�lɫ�H􇆑�����
e�1>(���L'0|���, ��J�����3��ٞ.y@��k�	C���3�BR���T5��(���
��Zr��� ��&��9�4�+X�.��N��g��% SZǩ���LrGI�V~N��N���W�V�yk�(�Tq����ۈ����iS�y5"'s��	q0nd�\��z�@�������'�K+UT@���T!a�s��[G���ь��@?\-�Ņ\�ŀ�:7�Cy:v����<�`s|LȬ��2��2��mG�{p��v�	��O}Ag��:�hI)� x-q/�6���$��5; ���'�ִ��f�n`l��If��#�cs[�����j�� �P\(�pk9��߰��� 3\�q%+{E���Q�'=���ml-p²(:�1~>�����]$bK���*�(��X�c�Y���K��8ny�)��  ���t�,�����ir�.��@�Uhw���/\o6����L���qG`h��(�~���A�F�b�)��Λ�v����Y�v�1� ��{��VV�Nb�Tc���V&�ݬ}��@uz�{{>��R�b�Q/ӃZ\�����l��{A�wbL3Э�o��)uTB����j�D|��C��_��SE��	��d؜�"�'Z0I��"y�Hm91c�-{�25�q�r�.�$��!�}�r"ٖ��Th���ꨀW�U�r���X�����j���ޓ�;k���<r��~(~ۉ�$�w0D�V1�nh�rl�d���ˍs��Kx��ِ��OaT9�-�s��arƬ�lKr*��)���#���/�l/@	g�X��Œq�a�!2CB5%�`ߡ����rk���ܒ��]����y�`���z�iJ���+����֙1l�4U�I66��mM�{ ����Y~�u�I�}��y�㐈�7���C�Jl �6~�+��~�ez�fR����1qN/���暈lko���Ը�����%[F���au�O��''=<�n��f"V�������3�씗$�`�q@��c�<B��#�Z �)��:���$�~�3L�E���b/�J�;A�܅��)�v����[�'g+]���F\W[�%�b�`�4�[��dr�?�o|*F r�� �"���X���l�kyH��"� ��y����p�%n�d?Y�q��!^i�{l��C���n�~���z������8]:�1_!�a�����.t�-�6y=l&T�j�pjx4E��f g�ܯM|�����u�$�gL�e�B����`-[}q4�$p �:�=���覒:劝P]	�H��[v��n��C�"�� 9|@�Y;|b��~��v�%���%�ļ�鲅0bO�2�j(���Q^H�%B��b�h8����-p:�a�mu(9�,�>P×��A��\W�g9���H�DD��$�Y�S�&
%7�xc���H��<S��-��7�J<�3I�a��
�۠8�!�(aM���?!�]b�X'�$�︔;iF0?�0T�p�&H$h�	�1ɖ℉�24�l��vY�F�����h�d�#���>R��@�at��P�Y+o��yZ�:���ǵ�</̴m�]��	��X�ɡ]���w�v$6D�~���r���;k���C���J6ωLbt���A��et��=�����,o2�B�`����[��D�����IC|^Q8/1���A)�FQ�S�]��z�Q�W����W�J����l��#>r�3�|�5���2X��`(��ڽ9�o�2��O�^�� {A�xЍ������=D<��8nJ��Įu��K�g�j��ɮM~E�u�5!A9,�T�"�R�0��Ia��t�j��1{Z=A�qY�"�l�0*�>9ǌQ�`��0���Z�rS�q����ݷy�j��R>��<�Lv4�B�[�/�@�Y��k�����3�c.-S�`�/2� �.�v�+��0��֚'wYE�;5?�l����W;!=vc�I���]0��e��c���=��$}�z�R����f?B��{�����o1���2�{����y[u����x\�x}���zÙ�{��A��RBr��iJW���B%]G�M3dnwgc:�s-E��̒�?�Ʒ��^�����3)�QU,J�T��Ȧ�N�,$=�1�Y����#f�V�r_e����z�ڋ8x��2��
򩰦���u��
����f���MIxzBژ�d�&��6�ʢ�r��+G $න��6�D
}������4\�������1�Μ�?��ZIj��M -b,]=&	��U4݊��+s[��86��NB�^6�]�@��UK$���`�4Y2U�
b���X;�M��)@��_޷7��u�~w�N�SzAR(`�0�������;�r��.l�P�\G( R䐭	�C�%�����[TP�4vg�"q�(
�i�ie��|N�G
���M^_nN���p�Zj��4���������{��N��'�"��A��$*'C?�Ļ��pI!$,E�����óAb�8 /����9L\Jǩ�__�5.�	v�r~Mxx!'��SWZ�}�N����z�8��)�(�٢L��$��>��g$�y���9���%<V�T��\�Ⓚ����(����pD�!&�p��ӹ�|�M�`s�cc;�|���lz�cg ��:g����:��#(�,�]�3�kD�?%ݬ�a^/ף��_S�|����.5^�Ĺ�&j �/(T�g�W�z�r�RdwOG��֢4Z�1O,S�;�I,���)	�����) ��cK%�p��RZ�U��v�a�ar�Dj�M�5�sGlD�W�tq�c�n����RFUh��w'y���ݽ��,y�K
�}��U���2%��0KX�qc_"\i�V�D�3��O���O�����[�W7pV�|͸E�&���;�F�)�j�Id4���=����+��,����1VnH?]4SMH?���u�qY�Dcl�t))�G�Ѹg>�'"���ь��Sn=vv����k�Acu#�l$���v*tZ�ș>$";�oF{��a��P�s�X��Ֆ͒����u(d\��55��b�m�d���Å[:��|g��|y4��x6Z4��M�-�	Z{
�]��3��_]�4�ȴ��D(�stƁOUy��(}�dҕ�BO����gp��#����x�|�D�/
�%���RcLRM'���6�p���|k�x�bU��L��d�b
⏁ ���4��O*}r������W;p���9�S��4W�!�zZ�`�k`�.i��Z����	w�C[K�v��T�$�Z|~��oM�d�}_qF���d���᯿�sO=iJ�$�*X��������6������m�^�~rFF08F����h)��"<M��U�ɪdB���C���^}}�ٟAFg�4j�q�1��F����1U���$U͢Q5�mfL� bc��M��MY[��T�\OZ�C�+f��pY�n��Ў��|��k�^���cIөA����x��3`z��o�B�L��Q �J7 �F�=�\B�2�@l'ϴ��~h�7���
g���=Ȭ�.�7-s�p��;	z��6�y�q콟�Q�Sc�u�+�8�i�SN��=�JQvNղ�9�f\��e�dd�hS�������P/��C�4zuq,Ek��ih�\1A�t�:؎245���-V�z ՂK�K_ʧ�H�2n������K��?����=b~�*,��%1����Ea��= �F���{n��:�	X�PfP�Kr-����"��E�F_�͞r=���o%UWp�6�O��}HO���d|��-s��`�2U{A/Ԫ��
�c�Z��nr�f�Uə�<��ED�����������-⢯}!ݴ(;گ��v��&.Ϯ��`�M���Q}rX��lmN �^I��`V#S�PG�X��HV��>�}�~ĸa��
��X���@���8�h�7s��{k�j�D�ܬv��:���M�*��W+|����aאjF��=sO���Ƒ���*����߃N� �4��&�o���jGҸ�Yl�PX*�yU�ܢ\~���X�.Pt��K�"��Wv`;� V|��Z�2~A���ű��2�L�ɂl��I��Ż�d�7�4 �x��J���'9�[t�,�l�֯h�B7*�9Y�^�ӳ�����Pˏ�
�	.l�Y(��f��X��g^PT�%��ۡ���#!س	���TEL��Z;�9"uz�@���{)Lb?�kj	P�b��1ζ^�߬�x�!b�l�w�:�y�c����X�@
�wp*O��%�.����6��U�ICQ�!Hܞ�S���ruD�kx�T~��?���cd�J�&y�K%���~���k�`n�`GQ���=�$/�lJuP_�,� ����ӀbL��s�!�G��a��od�3$������IH�����G��ѓ��䪙|B5�H�^ F2�3�r8�u��Ū�N���l%d�}2a��r�D��3��q�9�>p'e��g�>��k�ؾ槹�&��R�� �xx�w�˙L�)���2ºF���k]�n �}��`A��P�V�=(��2��C�K�$��'���u�qg�J�d�1S�{��<��c�E�m)�e	�w1�g�g��ҹ-�v���#��U� �V ������+������j�[�5��6&0T�hWh����Ĝ��(}IJ�rO�W�-�sH��a����HG�xf��o�