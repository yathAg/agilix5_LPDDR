	component ed_sim is
	end component ed_sim;

	u0 : component ed_sim
		;
