��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$��4�o;�����~>fF��i7����l`Û�%�l{t�r	�@Em�,�B=���Z�Vi�?�v��P�U�=�
��ۅf����u��ɡJמ��+"9e)xpƱ�7���r�CƖĽ-�=fK��ٞ�yq|J���\���t��(�B�^�=�S���Ȝ��܊6'{�߯AI.a��`=uzmu��g\'x𺼕�͢�*�g[+�CwT'r���ӱ��*��[��B�g�d��׌w���G��2�ޚ���l���P�����sk���ц(t�e�~c�d�����������5��	)�"��X��IUy�����ڥ�(����:��i�R>�M h�}���.Q���@S�Wpk��i�j+���U!ȱ�yf�R����[g~�˵��U?y��i��΋E�Aؿ��rƢr�I�˳��4B�UP�x��<�,��/��&f XŻt.���q���O����9֬}Y�P��D���	�⧢�i�Rڨ1%R���JV��.s�oI (� ��}�DU��Ҩ(�j��*}���)X\�欹oF������a!�d�K}�� �AɆ�;��A��{���ߖ}�뽠s� �I�Ј��4���D�9C�]L�����Σ�[0��;v�=1��u�1�|C�����ITb��>���D͏�7bo[�*�w��k��|� �Gb*k\��l����Tb��=�:Kӽ!������>�w%�[��	��t�u�r����7ړ���u��kȺ#����O�?f-t�&��k.
�!oşF�})���	�jMB�T��gV��`@t�fK��'��4�H6\�h�z��@�^2Y�NĲ'%�|�<� Ϲں��:����<
��4�V��LWd�^�8p�LJ��X���WJKP7Tj�ܲ���.V���"��$�����Vt<��F��q��֘�S���Z��]� Yz^H$�`Z�F|~�]��agp���O����H�r��0�jZ�)�{�^��f�	�7I8��g��u��^�����2p("�4���<V�~�|R��@���*n�-��6Sj����ZQdCEז��t�rC��6�\��+/����-��	��I���7��u:����ߟ��ޣ��0���3�G��>=���,��NY�GaBlF�*֮�:�~$yq3\����}���u?#��ݝOG%����yf�B��-ʙ��+��S��ퟹ鬶��-�n�3\�Sz�H��� d;�ݐ�â�a�Ԃ�:V��z.��O?����	��0���sj�2�A,��c�/�W}�-Q���]� ���7�$ܦH��R��Q�]!�����ji/�Q�� �,�ߢ��>^xnA����r$v`&ޮ<�)���\�,���?T��ʎч��E����@��u{��͋a5C�*nG+�ߛ���^��:c��u�Z�e�g�&bcʧ;�����_�q�r�D�݇McO���4�k��]�XP�M��ֈ|�%o*���H[c9/{U4�,���	ɘ��)��J��E���X>,^�,[�	��e�9��_�Я�Ž3�����엋7�]h�|� �;:H����]��[���F>��U����'�VD��R�Z�L��r��G�*�a��&}��6�?�0����b��7n*7����9y�K�r���KC%r@�DL�!Vm�((�qD8c�������N�j�%�{��ua뱠��/�VS:���B\�R9���饶���}�s?v�֣��ư�vz����<�δ���"3����Tƥ��r;��C��(6{ fϾ���'Q��6>�ؿ�!��G�ٜ���L�~-�0E[c��A�F�S,�e��W<����Tw��V&Y�᧑$�]�o�֥oۘ	��H�{�?\��0c�TLU ��ݲLj��mY�ѩsȕ��`c�c��mw�}���GY���U�Y��X�w)��&��k��pm-�U����ST\ӆOrv?<lm��E
4 �5��?n�6PѾS_�������$M|E�4��j3rƖ�T�Y�u2�dt��m,��S�>�/$FȽy"/t���� ���	l����G �J��c#ӹ�#�l�e�?L@��߽t��cj�$Q������˒%R��eU��r�	�v�ܼۛ�^��ĕu>a�����4���=zA�Lx�Q�q�1Z�*<�=r%���������fo0��פ��_�A�8D��BOֶ��&�T� Jg�iry9�~s�w��>�FVr� qy��X$��g��z�E(�V������?�7��$�U�]�T�8Las Q0Ɓ���9����j�s��f{ٻ��0�-�`�L(�0�|��q��3�O0����^m�K���Uؗ��
���x�FH����ɐj�}���(��_���T���F�r��7>��rJu�A}�����F�J1<��Û��`���,����u�D������ŗ˨���I���sʸ��i�,�Y��PL�X8�,�`T�r�2ߣ1v�������x{�Բ��o���nɉ�t.K�c�	��w�\GV�҈�i���#�z��x�w��`�?AQ컉����EȤ��O	V,��1∜�p�^܏��9.��[����ɺ�e%Ъ���7��4��)e
XQL����6����)����E�<k��@W�{$)���JLI\U��P��p��-�XH�3���T���N:�Y[YAu�g�!cGyӅ�3m�I*&�q5���]U�ӈT˚����Kgi���r�7�c�X��;�VP%�U��z�`�w�I��PQ����9b��y�Y�� o?�N���|�9gyEiv{�b� hK�c��[|���uSl@1!d��T�R�dJ��Cc�������]K�*�ϰ�-i�pZ�^���HV�4�t�r蝋'[�_����GS�r2���F>'�N���X����}���Ԣ��U�C��������Ժݨ�m�k�j?h2[&9w��^�����m��Y�e�*3ʺ��ǑӲ�����8N���P�(=A�46�ݗq��A�⁜�ܘ�]0�(� �}��l�s�n�"�����vZ���:^�+���k�0	m��cgu@E����,f}7V~�I��Q ��	[w��f���1�,HvK^��U�5�6�?�C�1(�B� ����6�Ҹ��b��v��I�f�����o��C�oa�q���~?ڏ��0t�{P�?	%�'+K���Ϸ;�|�cmC��O�Ԓ�?��"�p���|�Ӭ�<�8AW��f�5���Xr�,>(80V RJfZdA#L�A�&��E�G*3A
�i�F/��	Ռdp)M��zx�n�(I����I��PU��9ȋb4.4�v������S�c��]v]7�8�A��KN6!$\�T/��S���CG�	}����x��{yc�Ny�9Vsݱ[+�x�l6��hB�v���T���Yb�*�Țן���J��!d"d��`�c���r|~.������m��Zs���ՃG]v��R8\d~h��� n4��vD���$	��zB��*�8�m-Q�ˆ�g N��Xc���A`�@B��3��ׇ��Y��}9���E�r�*b�����%��;��/ȯ3FX����_;��H�g=�4s��v�����U��sCgŉ��y�Q�ۆ���ڗ� {P}*Ruc��RZoIK�{�L�i�_h�TQ�_3�].0�Nf1I��\8���[҂�nҀI(�-} Ԓ�@�Z�յ��X҉F��56�e\���y� <M��q�����9�V�i��21ν��������a�G�"���5 ��W�I��@(�@A�"��\����� �A,�Hȏ�JpY�Kb U;��E�>�1q8�MT��nw^]eh{4�f�T]'�y���������du<w�������?M:��༸gq�@ bx+�7ԏ*��$��V��3Y�կ����2�E��V
�EOo�]�c'A{���[�A�]�7��ת��M����4��7����1:�|�����";�M}�u����Z�^OXd+�r
9ޱ�?�R�w��d$���_{��ep/3���:�m1ws��`�`�,���E�{�D�f��d�F+�;`����Ժ��[��k?DD�+����A�W�Ƹ=$���]�2SI�Ծ��8
�ב�WY-��4Gk��ʍ,,�ݤ$��9������I��W��O��:�o3|P��v�𵔹���J�� �T�N�h�܇�o��ۗ�:T�\���W�Lɱ!ߟ�EG��˕��팖]�B�*�#"I��;�����~����`pX��	��<r��z�]`c�Մ����,;����
�
��4����V�9��w� {W��G.�"��'X�ig�`���NP�m\�P,z\m~]�[�4�2*Wx��d�
8h9��\I��t`���ml��_� %R8�����Pl٘��ò��?�iuKE9p�-�/��e�4l8�4�v�3
�l�vʪ|y`WK�ӲF�PA _@0�O#&�c)0�P�[��=��ϭ�>A�j�$��A��.�{�n����XxnC�}�D%��e�^:�YxN5� C1!�b�^|��o����{�8�%'�qi�g�R��Jh�#��g:�)`"%�e���5�%I���K``�X���7s�	�&��͐.���?w^��忛7�;�D�Յ���g(���{��������`'Cf�
*�>�K~^"���u��LtԞ�e�lJЍh�3�v`h;{.$��W:ֺ��-#���,WpU�W����/�!b��Y�􉒽/�O1|!�M,���e��({�q=9�RtM�+_Y2���&뼤!Һ�ᭁ�wQ�Tl�ok?'��C^�ud�<�B�Y�:q�&}r�
��粐E��TL�Ecs�w��I5ԅy���J���!|�2;����㷴�RW�K�I/x�8���\\1����'6bl�
�#i���X��a��Ӱ�J'EQ�.U���q��IO5�Kc(h}Ә�D]�S�#}��0��	��ը��b��yw�5v��ŭ��^Q�a�9�W_[')0�*�`�)b2 p��{[���]��|�)�1 R3G����e� �T���NA
ޯN)��/��`�����ͽu{���A�j��c~�2�)5�ܽ��H<�^�}X7������Ft�U�[�-4.�Y�ŷ���͏;�|�Iݚhtd�!l}l*��������B��/���M%t�HS�.{\|%�K�����+�S�X�*@#VE���<��W`�ΧY8$�y�H��E]�~"1�s���ù�}��
Q�;s�Ғ�|�	��~�%2��t��͋u�?��	[nX���L2��\����#>uW;c����yF"����h}c�)�_Z�A3��$ԓm���ajǨ!���3�ɽ����;K�J��O����W�/�>9ޚ7��fVV�z���Q�b�9�+zXt	J�������Tڇ�B��]����4�$�wC��Sy�5Zh���Y�ۇqʅ�a"���Z��h���p��,u�0��4a���uW��T���ߏ�E�%��u�J��B�[UrC�b,I������.q[��ՏvPOՂG:��X�_<��KS���f��m_�C�P��jY� @p�]j29&�� ��"��CVm<��rF;?wC\z�b{i틣��9��ih6 }x
��X'��J�o�Bg#��;F������0Ů�ּ�l��E�eX��vP�)�X�17\�Q��T��]en�>g� �5�p�|^Li3%���o��v�X?�G�Cؼ���l��-OF�����Rȱ:�P��
Ѝ�arb�"�j���^:�V+�i�I0)C}��IV��9I3V��=ԫ*4&M!��'���xf� �*�)�?S��<jv�E?�?���o��s9�Z�ܶ��pc�6����������ܴ�){�Oom���|dO9{�s#�-�1��K��h���9e2ܜN�ccdC��d&���J�,mƨ� {hx'j�fz!"��
�3u*D���^]�a�i�$�Pޤ�3\'v�����{q/���¿<�1���[ZF�w5�V4��r4�^�L�:`5���H�˘��.�)��]Y�'�w�'	(sE��s�ȵYkn� ��7ܑ��,'���B��������+<F��"H_�}�Ȗn�9i3�c��aҏ,3�5��Ә0:�[OE'�yq�0�}��_�D�{O�&��-r��|�@~i�H����L���/Q�#�u�3H����Z�� mQt�\~%V!��T���ɟ�&M�i��YN��,�����y��ǵ*�"��&2m�9/#�%�wlV�6w��������Ϳ���
ၸJ%1� �h:bM_V?�{A����Ʊ�@�&�|t祫FC�J�3 ���C_ODNz�0�$6?]�E�>����F��/V#[˄M����m�E��xխ�Xb�q�Iw�>��Ә�]��|G5bQ�����x�C�
���� �������4��+V�Sݚ�[����6�i�|��!�0� ��� f?Ǣ������l�ß�M�
3�b�0Q�`��.����sې��$|���NMOY�mɬ��	�M��Z�+�=��'Mx��!
%�����0/��yWk��̾;��y.��j�)�4%$pV���t�`��E��ܦ ���hX�Ӫq��@�p�c�R�c��mډ�� �#Hl;c�u!�z+ �l(��Q
�B�i�����@7N���}K-�O:IW3+��$�h�C�Lw_�?��#��!`��ߑn�ao#�������n��ݥ�ʕc˴�N��� �Yn�t�6��T��I9!��Q�-Ik�� �~UK����`8d~jA��q��ģ)wb5q8�"Mv��c�Fj%�����1n��?Q}�h<;�3oQu��UjC�D�F>g�	/A/[��I��XȏME��夢!�u��m�uf��[$H)�����2�?{&�Fs+���Wz��IZ�ܜEs/�]�)���^��@�R�x_���m��Ww�{)CYEDfz �Q��]�&�K D��!+�wW�zAp��N9)Ԙth��]:�c Na��}	0�w�[�<Eg-Qr��qL=��]A�P������<���ֲ��K���g�?l�xΡLo[i|�B���G�gc>N#�T��+Χ�h�R�oHJ�蒃o[1��j�;h[�]��9�(_��$A�h�z���s���o I�d=ϒ0���F<J���{G�e��8rJ�� �qt!������cD�y�7{_��a��Q�R��i��sZy���d��0�J-h��
c��s(TX���DA\+*c(P�z�B|ʙg4
F�{��q���R���n�Ƃ�g)�l�C�l�n�Σ�4D{���I�Ӵ�����Ζn<sf_� �k�)w��Ua�<v���3�v�CA#�DH ̙���$�]��0�I�1?K��3�a�%x�E�}zdY��>��!�.�]�ڰ�8��Y�F�IM��I��:7�n(1�M���6&��(���bɓ���F��Z��Q
a���c��u�	��s�E��P�+ݭ�xQ�Gȓ��??����rʽQ�d�
�����L:�mN=�h�}�����f�n2�o�qx����_�Y�)�������!�?�8�7���;x�W���{v�g���S�����L��	@-�<O���6+;���]$�lz���6�d�r��"�k�Nۛ� �H)L���dc��tO�ˋ"��'����������#����:��������;0f��k�(3�Hde�A�,j
9���&j�练=�<��_׷V���4�<��#cUDo��*T~��4PАX���fjn�2ڧ5cf�c�;q�jp�;�����dR��c,��J*o@p�|�����"��Yb!���5��io>�Gc�	ɍ���$.<�$[��6�*���1���aY9*�Nf�_��%�b<��H ���z���cvkp'�%3FvZ��A�Ou���B	�z9�A#+=-���9勼���8�W��u�wdڡZ2Ί���⯏y�1ƶ>0�]�IIp�じͼ�j�)�M�y�	��j5��6H�2�4c�� s٭c9v���ӧh��)�f�K=�B��5B�,�f5�n�|MS�t�GT�l�)i�`LN������`B���kQ@��HuBa�̘p�D�������H�[Y:=�˪��aDLH^i�#'����֨�3�S�*�$��a�����l���`VG��)�*꯲�k-k�
	>�L��!���'��c�RLߊ�Q��P���p�+��V/X*� 5���lB<��9��a�'�6`���d�{�"�Ѣ��S��(��]�q��F;Yi�˫"��y[(}�!J;���,�Bx������+�j���"�yPv�g��g����U�dN9�ԩ]�k�?��@��}(O�m���"�w�8W��<B�˚�G��	��� �iVk��3D�q���ܝ��\���#Z� W��Bw�:�Jt�̲�e��*�;���j9֝*���/�{�"Sr?�d�%�*|	�jЃ<HZ�@V�t�k�����3;#�m�.���Ę�.�)s�eFW���%Z����/����At>�-àJI�vͦnOt
|�Yӕ���!4�[�`�(^��/a�� a�c�ފ��!� �z��4+��b�Y8��Q?����@���|���� g�`�۾r ���}�б�U�BH֚�����RA��?&
-I�!oޏ�+��;wLM��l����=�<ڜ����X�FX�Uk�(F����&����4n���{q�u�޾گ�O�ۓ�y�� ػ�)��P�MIR�j�Z^�(ˑ�dc?��y�� s׷���7�󄋁�Cc��Y�F)����+�έ3jw��K��,]��C����n�[�k�R}'�x��?<Qm˳ar���e"��'��`�T�f/Dh��	��\�&�X�	X�%n�|���i%$��\�s���X�}��iھOk��:hV��~S]j��Y�a�v�̖�mu���$�=t|g�$V�\������9�`���`q_tgp/�������j���fO������#���S=κ���k�"�85���p�,����W�-e�mN �i0T�c�W+:���^�齔�I���7}1Գ��;�{r|�������2��A9S�*�=��G�k��`��/���B��c��mM��}'�˘=����(-�/��Pz �!�����d� �X�j��!hs���o�6\I�U$����ҧ�0�޹�qz@J�Z̥��5ÅC��|0�`�V�-7��2I���W�$k�J������`��Jb�z&����>�M��yR'�.���@�X�B�J��� ��`�g�ȶ:!řfݣi�=��j Kb��k��bJP�BO"M��*כ�~�@k��/޷>W�Ul^xv�v���I�>�` �����;� !1�'x�_^���Ŋ@����p�� F�6i��q�����/��ۇ��@�jO�i� ����ǜ`�[��1Z\�m��ʸ�x��޸ߨ��_��o�b%������¸ߕ��'�yn2�`�$U�������TF���%P�Om�b1peO?�}���t��W�S���i#ʤ �AkMZpS���Gժ%۝|��3�˙P�}�y���X�9~_�v+w|���9y1�o�HrV^�"@��ED}*~@J�^#{k�x��Vo���)��`4\/ϘVY��3�&z���`��8ԜVc�,y1��!^dJ@�5��3����A=�~j��`Vd�^�&�Q��N%J���MGrA'��2:�"I��Io�\D8�a_J���&!�LQ�)J�c�SG���<X_r;y�\	lB~�ߥ.e�S����ݰ �p������Ә��Q����X�.|��e�o�m)�[����
��x���*�^~W8�?�예�K�����j=���A.v�?��]��hJ���9"1a�_�r���Ү������t�47�M]�Nݯ4��t�[A`�O�z	 ý������[)��aw��z���}.m�9h��	���.��i��Y-!=��닠 d��J��ӳ�+s�j��e��k��7�>�k�^�ߧ]�]��^=���~}�}얦b�%7{�>%�J�K.x"( u�K��A����Xݣd,���L����bq��(=���,�����,�TN/�S��т.r�+@�n&����X�2��W��Cp1�MQ�|�B���IJ|3���)vM�,��c��o(�����J=����7�I��O�#�2�<Mjݕ��O���V�p���"����#n�o�> �#睫1�A���F0y��0ݾ�V��?-�(�wd�����2L�8G��[�N*�Z�Fn?��hq���lϳ�ΩoVo���(��)[��z�0�D �Ba������g���ˈ��0���|��p�;��;�\���t�uV��6W�Ʋ���������,��{��0�J W�|XR|�1n7哎 ��ec�O�ՠ�.O��"��ϣćA�u�v��QC_�����c��٘[�9�����(G@��|������� Y���&�Lv��v�9o�cg���>��[r��\:(�����q�t`;Tj�Ԑ�J�,NfE������O= ��.���a�m������Z�,SS�`Sꐱ�!�#�7��vT�5/��<t&