��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$��4�o;�����~>fF��i7����l`Û�%�l{t�r	�@Em�,�B=���Z�Vi�?�v��P�U�=�
��ۅf����u��ɡJמ��+"9e)xpƱ�7���r�CƖĽ-�=fK��ٞ�yq|J���\���t��(�B�^�=�S���Ȝ��܊6'{�߯AI.a��`=uzmu��g\'x𺼕�͢�*�g[+�CwT'r���ӱ��*��[��B�g�d��׌w���G��2�ޚ���l�h6O�������fE�8#�A�4��V���6N'�������`V����Q|Ɋ��%V�ZI]|�#M��gb8<N"�O9�	t�SM��\�Ǜ��"�1�^;����_WX�_2Ѳ�J�/��+G�1t���.u����e���o=��V�.������
�gC����\ꥥql������D�+-����a ��:К�ck"�@�9 D%1�8�@�����b�G�p=ˢ��j~jμ�W��L; �n��n���_�P*�C�Y�(��٩-�U��-�D��ۯD��H����;�4�9/(]{���{f[������#^������Pړ������I�����p�Fg^+���V�A�m��G"�~�U�p�O	+@N��U�(Ŏ5{�ZG�`Wg%NF`�P�N9�E+�##U^ �� ��1���k�l�t�\b1��P2?wz�/�������ꍦ��yF�*������
<�dGݧ#���g���lӮ<2;���ް4��B:��s���}��h���-mH1�e�S*��hP�
 �-�k�S:�d�k���Շl�
XlD���f#��"J��|?����*�i���%��͢?"^@�@*���5�r'��7��H�5�ܜ�#	�:=e�V�K��͑ ��҅��!cb�G�O5��h��|:#�u��-2����Q�a�trϢ�\r��3�\���z�y�9z�M:|�G���(>����f�r�1��S�Jƾo�U�9g�~�/�?���X	�#�w���"t�qz��z	&	��A�I�b��+H1�����׃6��Nh��n��)����7��U>"����S4Z'�7D&�u�E�*>��S�L��׊ٮuOq��%���{S����;��$�m����A�˄��j���ML��]���%*�v�o_�"�t�J
h�~��9��PI� � v*��<XM��~?v�`��bJbϡ6M p�Y���aj�B&�(�}x��`�3�cq�~䵥�!�_2A�E�N��2��ٻ�k�k�H�^�q���d���6�X�)��g����
U鷼�ᾥ�L���ȉ��ڂ�Q|���K~��	�(�'��W#�SK�� ^cd4V�����H�Bi��J��"���!5@�fSCd�uEl�$߻���s�6�u��(��X�y�W�tTh�O���/ì,*+��P��z�5#/l�y�PTO�'�,��h���R�Z�:��Ր�OMs'j"%����������W��������j���r9H���H�6��͝�8��)��mD�:CY�7�4��sLF0f���ݻ.7��"���)�p���)�lt��qb�n�2@�o�� �d+�m���!-�R�?��QNG�*�!��l�]j�m�����Th%i��S}�ΞXTVw��)���W(%A惖��+��J���)Rn���tt�S�;�`���@Xu챖0q���eQ����"]�f���PZ2J��L�o��y��1��>�r<c慷��� HL����n�b�<��Յ�M-&"4X�">FI��A��RТ���[��(�c���f��6��4=�5�Z$ry#�x*֖����~��Pš�$?������N<�wk���B��
��PI�9�dtv�׈+,� 5f
D�+����ۚ��Z���R��W�~%/qD� �p��7o}>�7&=(\ݵ��xZ�wA�<&F�f����	��,�a�
ް{|�ǚ��C�'u��a�4�G搒|ӓ�b�.V��*����Z�yd6fS����[�� ��Mޥ�b��������������38}�&s���B����i��:����ͅ�ΟЮj�\��r��R��sY�dYJ)k0g	���x@}5Wa�*�
r��=rs�PH��M7���}o�Q���� �r�-�YMi�-�T�0L�q�n����"����ǭ=V�t?��=(����.q�ѳ�y[�A�4!f� �k[���Lխ"�+���g�����%�i!�+�E�!zm�k�0�2��A�q�[H�2Kqڌ:�J�V�4����͟�/�m�Kt�4�2DC�m�/0���,ޏ@G�{��ѥ{µz��P	3f���vQPs��[j����㻣�FP��DpC�=�������n:�Pz��@֘��@���3���"<��K��3]z�l�kק�y(��ι���ek��M�^��?.x𔘲�K����znǜ��5n��57ߌ��XLW� .~נ�&\�
|�C��D��څ������.	bA�>(�����-�K��b�5����U�Y��k���n<yߖ�Bd�Q�03x����BE������b��4Zݯ��
���L��u,j��V�1�0�:+�ID��'��� ����&�>f.׾(	zb��#}�lߴn���N�,�̯ ���f��YubW1��l�*�;��P�,4~�T�O�����Ƨ&�j�5��n?	}QF�@�P��A �P�!7�܏��TD�������$�hk�(3W���E�Ӿ���-;����g��P��w� ?�٫����Z(\F>�4Y碇DW����uY��,�M��V4
�̺�p�'��?nTt������R�5�����,L_�_q�*�ǟދ��g7L}�v�0�3������Ǐ��q�q���A�/��q-T8��������|�J�"�=� Y�S<�E�*Ar%�W�%l��`P+�]�=ڲ��;�Z|�?�ϵh����5�,�q�Q6�(���@jB�X�E�P/�����NZm�2���Q�"t<7�o�=Q�I&υz�?�-����L߭9f����d�@ @��@���F��	qKJ]������hx�m�`�)������+bк^Þ^�W9MQ8L��H�m��$��G�Ԕ�/=�����v�b����JaحBR��텋3/oW���I�]mIj��ŗ���Ռ�y��d���|s�'�`��v�D!ś6�r���_�̋�:���l詨Ȕ)��{�n!\,+��/8�5NH/��:_��WK��+�MG��E]L��Z r���x���P~��3��-�9_b���.��I5���W+������R,O�Z��Q~6�Z��7�*o��v{��t��}�p��M�G��aگя[~�f/��P1�.v����j��dFY5�O�����s�e?��l��E��7��Z�ڸ�K���+��|Ѳ=�ۄ�B����1�&��=7���$��k?�a�z��p2�r�<u��d��9IK��b�n�HE������ �i-�2��O���\�@�I�`���� ?��`�4��fb���v���x�	n�"��5%2^�>R�{}�绺���H^4
�,�'ɷ��n��J5����#�(-\3�����3P��mS�v��39CG򫳗�Ѥ�Ѹ�,Ijdu�Z4�0m��\z�(X�m������Ӱ�Ɛ��B�{�3�|A�����)�u(S�*�h��^9��QJ+�+�ϩͷ4?�W�M�ֺ:H�Ϙ>���oM���7W���@B�)s�B����;���O��HEs��l&�Y��2n���K�([e�e_���td1�Ҁ�9[Ac��8�w��Ho��?k�5�,g�Z3�i{�T���:8�L�	�R�OSU��v�!�1E��4�똳����h"*2Ӧݭm;�]�by�8{�����~���R��'P�;�W#Zr�5�u�d
�'+n3���,�a���*)��/�w ��Lr���4/���'/�<�b������T�<=�y;2�o.HH
�lGs����|6ol~��s�kT��Đ�W�5�@{��_A�2E.M�ZQ_,R`����#�_�"E�V�wp��k�f}�gQ��v��D�wqx�N�(ۚԤ�Z�����B�%��Z�:ݪ[1 ʁN)z���¸���X�dg��}m_�}�u����~�]�p�핞S}z����������r�56*�5 x�s$+�㚨�A����l��gd梁�:$X�}�z߅YעMsAJ�����i��=��I�4����b}�eآ|?K�/v����6�]��~t �W'}��r����?��EPp��/�A�A���oNMq�vWr k}?�0�GiB"h<^X�1�UOo�27ᴓ���4�o՚7�^�8u�S���o�N���2}?���j��B��D�R��?5��_$��ey��!�(