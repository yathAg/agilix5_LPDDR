// ed_sim.v

// Generated using ACDS version 24.3.1 102

`timescale 1 ps / 1 ps
module ed_sim (
	);

	wire   [26:0] axil_driver_0_axil_driver_axi4_lite_awaddr;            // axil_driver_0:axil_driver_awaddr -> emif_io96b_lpddr4_0:s0_axi4lite_awaddr
	wire    [1:0] axil_driver_0_axil_driver_axi4_lite_bresp;             // emif_io96b_lpddr4_0:s0_axi4lite_bresp -> axil_driver_0:axil_driver_bresp
	wire          axil_driver_0_axil_driver_axi4_lite_arready;           // emif_io96b_lpddr4_0:s0_axi4lite_arready -> axil_driver_0:axil_driver_arready
	wire   [31:0] axil_driver_0_axil_driver_axi4_lite_rdata;             // emif_io96b_lpddr4_0:s0_axi4lite_rdata -> axil_driver_0:axil_driver_rdata
	wire    [3:0] axil_driver_0_axil_driver_axi4_lite_wstrb;             // axil_driver_0:axil_driver_wstrb -> emif_io96b_lpddr4_0:s0_axi4lite_wstrb
	wire          axil_driver_0_axil_driver_axi4_lite_wready;            // emif_io96b_lpddr4_0:s0_axi4lite_wready -> axil_driver_0:axil_driver_wready
	wire          axil_driver_0_axil_driver_axi4_lite_awready;           // emif_io96b_lpddr4_0:s0_axi4lite_awready -> axil_driver_0:axil_driver_awready
	wire          axil_driver_0_axil_driver_axi4_lite_rready;            // axil_driver_0:axil_driver_rready -> emif_io96b_lpddr4_0:s0_axi4lite_rready
	wire          axil_driver_0_axil_driver_axi4_lite_bready;            // axil_driver_0:axil_driver_bready -> emif_io96b_lpddr4_0:s0_axi4lite_bready
	wire          axil_driver_0_axil_driver_axi4_lite_wvalid;            // axil_driver_0:axil_driver_wvalid -> emif_io96b_lpddr4_0:s0_axi4lite_wvalid
	wire   [26:0] axil_driver_0_axil_driver_axi4_lite_araddr;            // axil_driver_0:axil_driver_araddr -> emif_io96b_lpddr4_0:s0_axi4lite_araddr
	wire    [1:0] axil_driver_0_axil_driver_axi4_lite_rresp;             // emif_io96b_lpddr4_0:s0_axi4lite_rresp -> axil_driver_0:axil_driver_rresp
	wire    [2:0] axil_driver_0_axil_driver_axi4_lite_arprot;            // axil_driver_0:axil_driver_arprot -> emif_io96b_lpddr4_0:s0_axi4lite_arprot
	wire   [31:0] axil_driver_0_axil_driver_axi4_lite_wdata;             // axil_driver_0:axil_driver_wdata -> emif_io96b_lpddr4_0:s0_axi4lite_wdata
	wire          axil_driver_0_axil_driver_axi4_lite_arvalid;           // axil_driver_0:axil_driver_arvalid -> emif_io96b_lpddr4_0:s0_axi4lite_arvalid
	wire    [2:0] axil_driver_0_axil_driver_axi4_lite_awprot;            // axil_driver_0:axil_driver_awprot -> emif_io96b_lpddr4_0:s0_axi4lite_awprot
	wire          axil_driver_0_axil_driver_axi4_lite_bvalid;            // emif_io96b_lpddr4_0:s0_axi4lite_bvalid -> axil_driver_0:axil_driver_bvalid
	wire          axil_driver_0_axil_driver_axi4_lite_awvalid;           // axil_driver_0:axil_driver_awvalid -> emif_io96b_lpddr4_0:s0_axi4lite_awvalid
	wire          axil_driver_0_axil_driver_axi4_lite_rvalid;            // emif_io96b_lpddr4_0:s0_axi4lite_rvalid -> axil_driver_0:axil_driver_rvalid
	wire          ref_clk_source_0_clk_clk;                              // ref_clk_source_0:clk -> emif_io96b_lpddr4_0:ref_clk
	wire          async_clk_source_clk_clk;                              // async_clk_source:clk -> user_pll:refclk
	wire          user_pll_outclk0_clk;                                  // user_pll:outclk_0 -> [emif_io96b_lpddr4_0:s0_axi4_clock_in, mm_interconnect_1:user_pll_outclk0_clk, reset_handler:clk, rst_controller_001:clk, rst_controller_002:clk, traffic_generator:driver0_clk]
	wire          user_pll_outclk1_clk;                                  // user_pll:outclk_1 -> [axil_driver_0:axil_driver_clk, emif_io96b_lpddr4_0:s0_axi4lite_clock, rst_controller:clk, traffic_generator:remote_intf_clk]
	wire          user_pll_locked_export;                                // user_pll:locked -> reset_handler:conduit_0
	wire    [3:0] emif_io96b_lpddr4_0_mem_0_mem_dqs_t;                   // [] -> [emif_io96b_lpddr4_0:mem_0_dqs_t, mem:mem_dqs_t_0]
	wire    [3:0] emif_io96b_lpddr4_0_mem_0_mem_dqs_c;                   // [] -> [emif_io96b_lpddr4_0:mem_0_dqs_c, mem:mem_dqs_c_0]
	wire   [31:0] emif_io96b_lpddr4_0_mem_0_mem_dq;                      // [] -> [emif_io96b_lpddr4_0:mem_0_dq, mem:mem_dq_0]
	wire    [0:0] emif_io96b_lpddr4_0_mem_0_mem_cs;                      // emif_io96b_lpddr4_0:mem_0_cs -> mem:mem_cs_0
	wire    [5:0] emif_io96b_lpddr4_0_mem_0_mem_ca;                      // emif_io96b_lpddr4_0:mem_0_ca -> mem:mem_ca_0
	wire    [3:0] emif_io96b_lpddr4_0_mem_0_mem_dmi;                     // [] -> [emif_io96b_lpddr4_0:mem_0_dmi, mem:mem_dmi_0]
	wire    [0:0] emif_io96b_lpddr4_0_mem_0_mem_cke;                     // emif_io96b_lpddr4_0:mem_0_cke -> mem:mem_cke_0
	wire    [0:0] emif_io96b_lpddr4_0_mem_ck_0_mem_ck_t;                 // emif_io96b_lpddr4_0:mem_0_ck_t -> mem:mem_ck_t_0
	wire    [0:0] emif_io96b_lpddr4_0_mem_ck_0_mem_ck_c;                 // emif_io96b_lpddr4_0:mem_0_ck_c -> mem:mem_ck_c_0
	wire          emif_io96b_lpddr4_0_mem_reset_n_mem_reset_n;           // emif_io96b_lpddr4_0:mem_0_reset_n -> mem:mem_reset_n_0
	wire          mem_oct_0_oct_rzqin;                                   // mem:oct_rzqin_0 -> emif_io96b_lpddr4_0:oct_rzqin_0
	wire          axil_driver_0_cal_done_rst_n_reset;                    // axil_driver_0:cal_done_rst_n -> [rst_controller_001:reset_in0, traffic_generator:driver0_reset_n]
	wire          rrip_ninit_done_reset;                                 // rrip:ninit_done -> [reset_handler:reset_n_0, user_pll:rst]
	wire          reset_handler_reset_n_out_reset;                       // reset_handler:reset_out_n -> [emif_io96b_lpddr4_0:core_init_n, rst_controller:reset_in0, traffic_generator:remote_intf_reset_n]
	wire    [1:0] traffic_generator_driver0_axi4_awburst;                // traffic_generator:driver0_axi4_awburst -> mm_interconnect_1:traffic_generator_driver0_axi4_awburst
	wire    [0:0] traffic_generator_driver0_axi4_awuser;                 // traffic_generator:driver0_axi4_awuser -> mm_interconnect_1:traffic_generator_driver0_axi4_awuser
	wire    [7:0] traffic_generator_driver0_axi4_arlen;                  // traffic_generator:driver0_axi4_arlen -> mm_interconnect_1:traffic_generator_driver0_axi4_arlen
	wire          traffic_generator_driver0_axi4_wready;                 // mm_interconnect_1:traffic_generator_driver0_axi4_wready -> traffic_generator:driver0_axi4_wready
	wire   [31:0] traffic_generator_driver0_axi4_wstrb;                  // traffic_generator:driver0_axi4_wstrb -> mm_interconnect_1:traffic_generator_driver0_axi4_wstrb
	wire    [6:0] traffic_generator_driver0_axi4_rid;                    // mm_interconnect_1:traffic_generator_driver0_axi4_rid -> traffic_generator:driver0_axi4_rid
	wire          traffic_generator_driver0_axi4_rready;                 // traffic_generator:driver0_axi4_rready -> mm_interconnect_1:traffic_generator_driver0_axi4_rready
	wire    [7:0] traffic_generator_driver0_axi4_awlen;                  // traffic_generator:driver0_axi4_awlen -> mm_interconnect_1:traffic_generator_driver0_axi4_awlen
	wire    [3:0] traffic_generator_driver0_axi4_arcache;                // traffic_generator:driver0_axi4_arcache -> mm_interconnect_1:traffic_generator_driver0_axi4_arcache
	wire   [31:0] traffic_generator_driver0_axi4_araddr;                 // traffic_generator:driver0_axi4_araddr -> mm_interconnect_1:traffic_generator_driver0_axi4_araddr
	wire          traffic_generator_driver0_axi4_wvalid;                 // traffic_generator:driver0_axi4_wvalid -> mm_interconnect_1:traffic_generator_driver0_axi4_wvalid
	wire    [2:0] traffic_generator_driver0_axi4_arprot;                 // traffic_generator:driver0_axi4_arprot -> mm_interconnect_1:traffic_generator_driver0_axi4_arprot
	wire    [2:0] traffic_generator_driver0_axi4_awprot;                 // traffic_generator:driver0_axi4_awprot -> mm_interconnect_1:traffic_generator_driver0_axi4_awprot
	wire          traffic_generator_driver0_axi4_arvalid;                // traffic_generator:driver0_axi4_arvalid -> mm_interconnect_1:traffic_generator_driver0_axi4_arvalid
	wire  [255:0] traffic_generator_driver0_axi4_wdata;                  // traffic_generator:driver0_axi4_wdata -> mm_interconnect_1:traffic_generator_driver0_axi4_wdata
	wire    [3:0] traffic_generator_driver0_axi4_awcache;                // traffic_generator:driver0_axi4_awcache -> mm_interconnect_1:traffic_generator_driver0_axi4_awcache
	wire    [6:0] traffic_generator_driver0_axi4_arid;                   // traffic_generator:driver0_axi4_arid -> mm_interconnect_1:traffic_generator_driver0_axi4_arid
	wire    [0:0] traffic_generator_driver0_axi4_arlock;                 // traffic_generator:driver0_axi4_arlock -> mm_interconnect_1:traffic_generator_driver0_axi4_arlock
	wire    [0:0] traffic_generator_driver0_axi4_awlock;                 // traffic_generator:driver0_axi4_awlock -> mm_interconnect_1:traffic_generator_driver0_axi4_awlock
	wire   [31:0] traffic_generator_driver0_axi4_awaddr;                 // traffic_generator:driver0_axi4_awaddr -> mm_interconnect_1:traffic_generator_driver0_axi4_awaddr
	wire          traffic_generator_driver0_axi4_arready;                // mm_interconnect_1:traffic_generator_driver0_axi4_arready -> traffic_generator:driver0_axi4_arready
	wire    [1:0] traffic_generator_driver0_axi4_bresp;                  // mm_interconnect_1:traffic_generator_driver0_axi4_bresp -> traffic_generator:driver0_axi4_bresp
	wire  [255:0] traffic_generator_driver0_axi4_rdata;                  // mm_interconnect_1:traffic_generator_driver0_axi4_rdata -> traffic_generator:driver0_axi4_rdata
	wire          traffic_generator_driver0_axi4_awready;                // mm_interconnect_1:traffic_generator_driver0_axi4_awready -> traffic_generator:driver0_axi4_awready
	wire    [1:0] traffic_generator_driver0_axi4_arburst;                // traffic_generator:driver0_axi4_arburst -> mm_interconnect_1:traffic_generator_driver0_axi4_arburst
	wire    [2:0] traffic_generator_driver0_axi4_arsize;                 // traffic_generator:driver0_axi4_arsize -> mm_interconnect_1:traffic_generator_driver0_axi4_arsize
	wire          traffic_generator_driver0_axi4_bready;                 // traffic_generator:driver0_axi4_bready -> mm_interconnect_1:traffic_generator_driver0_axi4_bready
	wire          traffic_generator_driver0_axi4_rlast;                  // mm_interconnect_1:traffic_generator_driver0_axi4_rlast -> traffic_generator:driver0_axi4_rlast
	wire          traffic_generator_driver0_axi4_wlast;                  // traffic_generator:driver0_axi4_wlast -> mm_interconnect_1:traffic_generator_driver0_axi4_wlast
	wire    [1:0] traffic_generator_driver0_axi4_rresp;                  // mm_interconnect_1:traffic_generator_driver0_axi4_rresp -> traffic_generator:driver0_axi4_rresp
	wire    [6:0] traffic_generator_driver0_axi4_awid;                   // traffic_generator:driver0_axi4_awid -> mm_interconnect_1:traffic_generator_driver0_axi4_awid
	wire    [6:0] traffic_generator_driver0_axi4_bid;                    // mm_interconnect_1:traffic_generator_driver0_axi4_bid -> traffic_generator:driver0_axi4_bid
	wire          traffic_generator_driver0_axi4_bvalid;                 // mm_interconnect_1:traffic_generator_driver0_axi4_bvalid -> traffic_generator:driver0_axi4_bvalid
	wire          traffic_generator_driver0_axi4_awvalid;                // traffic_generator:driver0_axi4_awvalid -> mm_interconnect_1:traffic_generator_driver0_axi4_awvalid
	wire    [2:0] traffic_generator_driver0_axi4_awsize;                 // traffic_generator:driver0_axi4_awsize -> mm_interconnect_1:traffic_generator_driver0_axi4_awsize
	wire    [0:0] traffic_generator_driver0_axi4_aruser;                 // traffic_generator:driver0_axi4_aruser -> mm_interconnect_1:traffic_generator_driver0_axi4_aruser
	wire          traffic_generator_driver0_axi4_rvalid;                 // mm_interconnect_1:traffic_generator_driver0_axi4_rvalid -> traffic_generator:driver0_axi4_rvalid
	wire   [31:0] mm_interconnect_1_emif_io96b_lpddr4_0_s0_axi4_ruser;   // emif_io96b_lpddr4_0:s0_axi4_ruser -> mm_interconnect_1:emif_io96b_lpddr4_0_s0_axi4_ruser
	wire   [31:0] mm_interconnect_1_emif_io96b_lpddr4_0_s0_axi4_wuser;   // mm_interconnect_1:emif_io96b_lpddr4_0_s0_axi4_wuser -> emif_io96b_lpddr4_0:s0_axi4_wuser
	wire    [1:0] mm_interconnect_1_emif_io96b_lpddr4_0_s0_axi4_awburst; // mm_interconnect_1:emif_io96b_lpddr4_0_s0_axi4_awburst -> emif_io96b_lpddr4_0:s0_axi4_awburst
	wire   [13:0] mm_interconnect_1_emif_io96b_lpddr4_0_s0_axi4_awuser;  // mm_interconnect_1:emif_io96b_lpddr4_0_s0_axi4_awuser -> emif_io96b_lpddr4_0:s0_axi4_awuser
	wire    [7:0] mm_interconnect_1_emif_io96b_lpddr4_0_s0_axi4_arlen;   // mm_interconnect_1:emif_io96b_lpddr4_0_s0_axi4_arlen -> emif_io96b_lpddr4_0:s0_axi4_arlen
	wire    [3:0] mm_interconnect_1_emif_io96b_lpddr4_0_s0_axi4_arqos;   // mm_interconnect_1:emif_io96b_lpddr4_0_s0_axi4_arqos -> emif_io96b_lpddr4_0:s0_axi4_arqos
	wire   [31:0] mm_interconnect_1_emif_io96b_lpddr4_0_s0_axi4_wstrb;   // mm_interconnect_1:emif_io96b_lpddr4_0_s0_axi4_wstrb -> emif_io96b_lpddr4_0:s0_axi4_wstrb
	wire          mm_interconnect_1_emif_io96b_lpddr4_0_s0_axi4_wready;  // emif_io96b_lpddr4_0:s0_axi4_wready -> mm_interconnect_1:emif_io96b_lpddr4_0_s0_axi4_wready
	wire    [6:0] mm_interconnect_1_emif_io96b_lpddr4_0_s0_axi4_rid;     // emif_io96b_lpddr4_0:s0_axi4_rid -> mm_interconnect_1:emif_io96b_lpddr4_0_s0_axi4_rid
	wire          mm_interconnect_1_emif_io96b_lpddr4_0_s0_axi4_rready;  // mm_interconnect_1:emif_io96b_lpddr4_0_s0_axi4_rready -> emif_io96b_lpddr4_0:s0_axi4_rready
	wire    [7:0] mm_interconnect_1_emif_io96b_lpddr4_0_s0_axi4_awlen;   // mm_interconnect_1:emif_io96b_lpddr4_0_s0_axi4_awlen -> emif_io96b_lpddr4_0:s0_axi4_awlen
	wire    [3:0] mm_interconnect_1_emif_io96b_lpddr4_0_s0_axi4_awqos;   // mm_interconnect_1:emif_io96b_lpddr4_0_s0_axi4_awqos -> emif_io96b_lpddr4_0:s0_axi4_awqos
	wire          mm_interconnect_1_emif_io96b_lpddr4_0_s0_axi4_wvalid;  // mm_interconnect_1:emif_io96b_lpddr4_0_s0_axi4_wvalid -> emif_io96b_lpddr4_0:s0_axi4_wvalid
	wire   [31:0] mm_interconnect_1_emif_io96b_lpddr4_0_s0_axi4_araddr;  // mm_interconnect_1:emif_io96b_lpddr4_0_s0_axi4_araddr -> emif_io96b_lpddr4_0:s0_axi4_araddr
	wire    [2:0] mm_interconnect_1_emif_io96b_lpddr4_0_s0_axi4_arprot;  // mm_interconnect_1:emif_io96b_lpddr4_0_s0_axi4_arprot -> emif_io96b_lpddr4_0:s0_axi4_arprot
	wire    [2:0] mm_interconnect_1_emif_io96b_lpddr4_0_s0_axi4_awprot;  // mm_interconnect_1:emif_io96b_lpddr4_0_s0_axi4_awprot -> emif_io96b_lpddr4_0:s0_axi4_awprot
	wire  [255:0] mm_interconnect_1_emif_io96b_lpddr4_0_s0_axi4_wdata;   // mm_interconnect_1:emif_io96b_lpddr4_0_s0_axi4_wdata -> emif_io96b_lpddr4_0:s0_axi4_wdata
	wire          mm_interconnect_1_emif_io96b_lpddr4_0_s0_axi4_arvalid; // mm_interconnect_1:emif_io96b_lpddr4_0_s0_axi4_arvalid -> emif_io96b_lpddr4_0:s0_axi4_arvalid
	wire    [6:0] mm_interconnect_1_emif_io96b_lpddr4_0_s0_axi4_arid;    // mm_interconnect_1:emif_io96b_lpddr4_0_s0_axi4_arid -> emif_io96b_lpddr4_0:s0_axi4_arid
	wire    [0:0] mm_interconnect_1_emif_io96b_lpddr4_0_s0_axi4_arlock;  // mm_interconnect_1:emif_io96b_lpddr4_0_s0_axi4_arlock -> emif_io96b_lpddr4_0:s0_axi4_arlock
	wire    [0:0] mm_interconnect_1_emif_io96b_lpddr4_0_s0_axi4_awlock;  // mm_interconnect_1:emif_io96b_lpddr4_0_s0_axi4_awlock -> emif_io96b_lpddr4_0:s0_axi4_awlock
	wire   [31:0] mm_interconnect_1_emif_io96b_lpddr4_0_s0_axi4_awaddr;  // mm_interconnect_1:emif_io96b_lpddr4_0_s0_axi4_awaddr -> emif_io96b_lpddr4_0:s0_axi4_awaddr
	wire    [1:0] mm_interconnect_1_emif_io96b_lpddr4_0_s0_axi4_bresp;   // emif_io96b_lpddr4_0:s0_axi4_bresp -> mm_interconnect_1:emif_io96b_lpddr4_0_s0_axi4_bresp
	wire          mm_interconnect_1_emif_io96b_lpddr4_0_s0_axi4_arready; // emif_io96b_lpddr4_0:s0_axi4_arready -> mm_interconnect_1:emif_io96b_lpddr4_0_s0_axi4_arready
	wire  [255:0] mm_interconnect_1_emif_io96b_lpddr4_0_s0_axi4_rdata;   // emif_io96b_lpddr4_0:s0_axi4_rdata -> mm_interconnect_1:emif_io96b_lpddr4_0_s0_axi4_rdata
	wire          mm_interconnect_1_emif_io96b_lpddr4_0_s0_axi4_awready; // emif_io96b_lpddr4_0:s0_axi4_awready -> mm_interconnect_1:emif_io96b_lpddr4_0_s0_axi4_awready
	wire    [1:0] mm_interconnect_1_emif_io96b_lpddr4_0_s0_axi4_arburst; // mm_interconnect_1:emif_io96b_lpddr4_0_s0_axi4_arburst -> emif_io96b_lpddr4_0:s0_axi4_arburst
	wire    [2:0] mm_interconnect_1_emif_io96b_lpddr4_0_s0_axi4_arsize;  // mm_interconnect_1:emif_io96b_lpddr4_0_s0_axi4_arsize -> emif_io96b_lpddr4_0:s0_axi4_arsize
	wire          mm_interconnect_1_emif_io96b_lpddr4_0_s0_axi4_bready;  // mm_interconnect_1:emif_io96b_lpddr4_0_s0_axi4_bready -> emif_io96b_lpddr4_0:s0_axi4_bready
	wire          mm_interconnect_1_emif_io96b_lpddr4_0_s0_axi4_rlast;   // emif_io96b_lpddr4_0:s0_axi4_rlast -> mm_interconnect_1:emif_io96b_lpddr4_0_s0_axi4_rlast
	wire          mm_interconnect_1_emif_io96b_lpddr4_0_s0_axi4_wlast;   // mm_interconnect_1:emif_io96b_lpddr4_0_s0_axi4_wlast -> emif_io96b_lpddr4_0:s0_axi4_wlast
	wire    [1:0] mm_interconnect_1_emif_io96b_lpddr4_0_s0_axi4_rresp;   // emif_io96b_lpddr4_0:s0_axi4_rresp -> mm_interconnect_1:emif_io96b_lpddr4_0_s0_axi4_rresp
	wire    [6:0] mm_interconnect_1_emif_io96b_lpddr4_0_s0_axi4_awid;    // mm_interconnect_1:emif_io96b_lpddr4_0_s0_axi4_awid -> emif_io96b_lpddr4_0:s0_axi4_awid
	wire    [6:0] mm_interconnect_1_emif_io96b_lpddr4_0_s0_axi4_bid;     // emif_io96b_lpddr4_0:s0_axi4_bid -> mm_interconnect_1:emif_io96b_lpddr4_0_s0_axi4_bid
	wire          mm_interconnect_1_emif_io96b_lpddr4_0_s0_axi4_bvalid;  // emif_io96b_lpddr4_0:s0_axi4_bvalid -> mm_interconnect_1:emif_io96b_lpddr4_0_s0_axi4_bvalid
	wire    [2:0] mm_interconnect_1_emif_io96b_lpddr4_0_s0_axi4_awsize;  // mm_interconnect_1:emif_io96b_lpddr4_0_s0_axi4_awsize -> emif_io96b_lpddr4_0:s0_axi4_awsize
	wire          mm_interconnect_1_emif_io96b_lpddr4_0_s0_axi4_awvalid; // mm_interconnect_1:emif_io96b_lpddr4_0_s0_axi4_awvalid -> emif_io96b_lpddr4_0:s0_axi4_awvalid
	wire   [13:0] mm_interconnect_1_emif_io96b_lpddr4_0_s0_axi4_aruser;  // mm_interconnect_1:emif_io96b_lpddr4_0_s0_axi4_aruser -> emif_io96b_lpddr4_0:s0_axi4_aruser
	wire          mm_interconnect_1_emif_io96b_lpddr4_0_s0_axi4_rvalid;  // emif_io96b_lpddr4_0:s0_axi4_rvalid -> mm_interconnect_1:emif_io96b_lpddr4_0_s0_axi4_rvalid
	wire          rst_controller_reset_out_reset;                        // rst_controller:reset_out -> [axil_driver_0:axil_driver_rst_n, emif_io96b_lpddr4_0:s0_axi4lite_reset_n]
	wire          rst_controller_001_reset_out_reset;                    // rst_controller_001:reset_out -> mm_interconnect_1:traffic_generator_driver0_axi4_translator_clk_reset_reset_bridge_in_reset_reset
	wire          rst_controller_002_reset_out_reset;                    // rst_controller_002:reset_out -> mm_interconnect_1:emif_io96b_lpddr4_0_s0_axi4_translator_clk_reset_reset_bridge_in_reset_reset
	wire          emif_io96b_lpddr4_0_s0_axi4_ctrl_ready_reset;          // emif_io96b_lpddr4_0:s0_axi4_reset_n -> rst_controller_002:reset_in0

	ed_sim_async_clk_source async_clk_source (
		.clk (async_clk_source_clk_clk)  //  output,  width = 1, clk.clk
	);

	ed_sim_axil_driver_0 axil_driver_0 (
		.axil_driver_clk     (user_pll_outclk1_clk),                        //   input,   width = 1,       axil_driver_clk.clk
		.axil_driver_rst_n   (~rst_controller_reset_out_reset),             //   input,   width = 1,     axil_driver_rst_n.reset_n
		.axil_driver_awaddr  (axil_driver_0_axil_driver_axi4_lite_awaddr),  //  output,  width = 27, axil_driver_axi4_lite.awaddr
		.axil_driver_awvalid (axil_driver_0_axil_driver_axi4_lite_awvalid), //  output,   width = 1,                      .awvalid
		.axil_driver_awready (axil_driver_0_axil_driver_axi4_lite_awready), //   input,   width = 1,                      .awready
		.axil_driver_wdata   (axil_driver_0_axil_driver_axi4_lite_wdata),   //  output,  width = 32,                      .wdata
		.axil_driver_wstrb   (axil_driver_0_axil_driver_axi4_lite_wstrb),   //  output,   width = 4,                      .wstrb
		.axil_driver_wvalid  (axil_driver_0_axil_driver_axi4_lite_wvalid),  //  output,   width = 1,                      .wvalid
		.axil_driver_wready  (axil_driver_0_axil_driver_axi4_lite_wready),  //   input,   width = 1,                      .wready
		.axil_driver_bresp   (axil_driver_0_axil_driver_axi4_lite_bresp),   //   input,   width = 2,                      .bresp
		.axil_driver_bvalid  (axil_driver_0_axil_driver_axi4_lite_bvalid),  //   input,   width = 1,                      .bvalid
		.axil_driver_bready  (axil_driver_0_axil_driver_axi4_lite_bready),  //  output,   width = 1,                      .bready
		.axil_driver_araddr  (axil_driver_0_axil_driver_axi4_lite_araddr),  //  output,  width = 27,                      .araddr
		.axil_driver_arvalid (axil_driver_0_axil_driver_axi4_lite_arvalid), //  output,   width = 1,                      .arvalid
		.axil_driver_arready (axil_driver_0_axil_driver_axi4_lite_arready), //   input,   width = 1,                      .arready
		.axil_driver_rdata   (axil_driver_0_axil_driver_axi4_lite_rdata),   //   input,  width = 32,                      .rdata
		.axil_driver_rresp   (axil_driver_0_axil_driver_axi4_lite_rresp),   //   input,   width = 2,                      .rresp
		.axil_driver_rvalid  (axil_driver_0_axil_driver_axi4_lite_rvalid),  //   input,   width = 1,                      .rvalid
		.axil_driver_rready  (axil_driver_0_axil_driver_axi4_lite_rready),  //  output,   width = 1,                      .rready
		.axil_driver_awprot  (axil_driver_0_axil_driver_axi4_lite_awprot),  //  output,   width = 3,                      .awprot
		.axil_driver_arprot  (axil_driver_0_axil_driver_axi4_lite_arprot),  //  output,   width = 3,                      .arprot
		.cal_done_rst_n      (axil_driver_0_cal_done_rst_n_reset)           //  output,   width = 1,        cal_done_rst_n.reset_n
	);

	ed_sim_emif_io96b_lpddr4_0 emif_io96b_lpddr4_0 (
		.s0_axi4_clock_in    (user_pll_outclk0_clk),                                  //   input,    width = 1,    s0_axi4_clock_in.clk
		.core_init_n         (reset_handler_reset_n_out_reset),                       //   input,    width = 1,         core_init_n.reset_n
		.s0_axi4_reset_n     (emif_io96b_lpddr4_0_s0_axi4_ctrl_ready_reset),          //  output,    width = 1,  s0_axi4_ctrl_ready.reset_n
		.s0_axi4_awaddr      (mm_interconnect_1_emif_io96b_lpddr4_0_s0_axi4_awaddr),  //   input,   width = 32,             s0_axi4.awaddr
		.s0_axi4_awburst     (mm_interconnect_1_emif_io96b_lpddr4_0_s0_axi4_awburst), //   input,    width = 2,                    .awburst
		.s0_axi4_awid        (mm_interconnect_1_emif_io96b_lpddr4_0_s0_axi4_awid),    //   input,    width = 7,                    .awid
		.s0_axi4_awlen       (mm_interconnect_1_emif_io96b_lpddr4_0_s0_axi4_awlen),   //   input,    width = 8,                    .awlen
		.s0_axi4_awlock      (mm_interconnect_1_emif_io96b_lpddr4_0_s0_axi4_awlock),  //   input,    width = 1,                    .awlock
		.s0_axi4_awqos       (mm_interconnect_1_emif_io96b_lpddr4_0_s0_axi4_awqos),   //   input,    width = 4,                    .awqos
		.s0_axi4_awsize      (mm_interconnect_1_emif_io96b_lpddr4_0_s0_axi4_awsize),  //   input,    width = 3,                    .awsize
		.s0_axi4_awvalid     (mm_interconnect_1_emif_io96b_lpddr4_0_s0_axi4_awvalid), //   input,    width = 1,                    .awvalid
		.s0_axi4_awuser      (mm_interconnect_1_emif_io96b_lpddr4_0_s0_axi4_awuser),  //   input,   width = 14,                    .awuser
		.s0_axi4_awprot      (mm_interconnect_1_emif_io96b_lpddr4_0_s0_axi4_awprot),  //   input,    width = 3,                    .awprot
		.s0_axi4_awready     (mm_interconnect_1_emif_io96b_lpddr4_0_s0_axi4_awready), //  output,    width = 1,                    .awready
		.s0_axi4_araddr      (mm_interconnect_1_emif_io96b_lpddr4_0_s0_axi4_araddr),  //   input,   width = 32,                    .araddr
		.s0_axi4_arburst     (mm_interconnect_1_emif_io96b_lpddr4_0_s0_axi4_arburst), //   input,    width = 2,                    .arburst
		.s0_axi4_arid        (mm_interconnect_1_emif_io96b_lpddr4_0_s0_axi4_arid),    //   input,    width = 7,                    .arid
		.s0_axi4_arlen       (mm_interconnect_1_emif_io96b_lpddr4_0_s0_axi4_arlen),   //   input,    width = 8,                    .arlen
		.s0_axi4_arlock      (mm_interconnect_1_emif_io96b_lpddr4_0_s0_axi4_arlock),  //   input,    width = 1,                    .arlock
		.s0_axi4_arqos       (mm_interconnect_1_emif_io96b_lpddr4_0_s0_axi4_arqos),   //   input,    width = 4,                    .arqos
		.s0_axi4_arsize      (mm_interconnect_1_emif_io96b_lpddr4_0_s0_axi4_arsize),  //   input,    width = 3,                    .arsize
		.s0_axi4_arvalid     (mm_interconnect_1_emif_io96b_lpddr4_0_s0_axi4_arvalid), //   input,    width = 1,                    .arvalid
		.s0_axi4_aruser      (mm_interconnect_1_emif_io96b_lpddr4_0_s0_axi4_aruser),  //   input,   width = 14,                    .aruser
		.s0_axi4_arprot      (mm_interconnect_1_emif_io96b_lpddr4_0_s0_axi4_arprot),  //   input,    width = 3,                    .arprot
		.s0_axi4_arready     (mm_interconnect_1_emif_io96b_lpddr4_0_s0_axi4_arready), //  output,    width = 1,                    .arready
		.s0_axi4_wdata       (mm_interconnect_1_emif_io96b_lpddr4_0_s0_axi4_wdata),   //   input,  width = 256,                    .wdata
		.s0_axi4_wstrb       (mm_interconnect_1_emif_io96b_lpddr4_0_s0_axi4_wstrb),   //   input,   width = 32,                    .wstrb
		.s0_axi4_wlast       (mm_interconnect_1_emif_io96b_lpddr4_0_s0_axi4_wlast),   //   input,    width = 1,                    .wlast
		.s0_axi4_wvalid      (mm_interconnect_1_emif_io96b_lpddr4_0_s0_axi4_wvalid),  //   input,    width = 1,                    .wvalid
		.s0_axi4_wuser       (mm_interconnect_1_emif_io96b_lpddr4_0_s0_axi4_wuser),   //   input,   width = 32,                    .wuser
		.s0_axi4_wready      (mm_interconnect_1_emif_io96b_lpddr4_0_s0_axi4_wready),  //  output,    width = 1,                    .wready
		.s0_axi4_bready      (mm_interconnect_1_emif_io96b_lpddr4_0_s0_axi4_bready),  //   input,    width = 1,                    .bready
		.s0_axi4_bid         (mm_interconnect_1_emif_io96b_lpddr4_0_s0_axi4_bid),     //  output,    width = 7,                    .bid
		.s0_axi4_bresp       (mm_interconnect_1_emif_io96b_lpddr4_0_s0_axi4_bresp),   //  output,    width = 2,                    .bresp
		.s0_axi4_bvalid      (mm_interconnect_1_emif_io96b_lpddr4_0_s0_axi4_bvalid),  //  output,    width = 1,                    .bvalid
		.s0_axi4_rready      (mm_interconnect_1_emif_io96b_lpddr4_0_s0_axi4_rready),  //   input,    width = 1,                    .rready
		.s0_axi4_ruser       (mm_interconnect_1_emif_io96b_lpddr4_0_s0_axi4_ruser),   //  output,   width = 32,                    .ruser
		.s0_axi4_rdata       (mm_interconnect_1_emif_io96b_lpddr4_0_s0_axi4_rdata),   //  output,  width = 256,                    .rdata
		.s0_axi4_rid         (mm_interconnect_1_emif_io96b_lpddr4_0_s0_axi4_rid),     //  output,    width = 7,                    .rid
		.s0_axi4_rlast       (mm_interconnect_1_emif_io96b_lpddr4_0_s0_axi4_rlast),   //  output,    width = 1,                    .rlast
		.s0_axi4_rresp       (mm_interconnect_1_emif_io96b_lpddr4_0_s0_axi4_rresp),   //  output,    width = 2,                    .rresp
		.s0_axi4_rvalid      (mm_interconnect_1_emif_io96b_lpddr4_0_s0_axi4_rvalid),  //  output,    width = 1,                    .rvalid
		.s0_axi4lite_clock   (user_pll_outclk1_clk),                                  //   input,    width = 1,   s0_axi4lite_clock.clk
		.s0_axi4lite_reset_n (~rst_controller_reset_out_reset),                       //   input,    width = 1, s0_axi4lite_reset_n.reset_n
		.s0_axi4lite_awaddr  (axil_driver_0_axil_driver_axi4_lite_awaddr),            //   input,   width = 27,         s0_axi4lite.awaddr
		.s0_axi4lite_awprot  (axil_driver_0_axil_driver_axi4_lite_awprot),            //   input,    width = 3,                    .awprot
		.s0_axi4lite_awvalid (axil_driver_0_axil_driver_axi4_lite_awvalid),           //   input,    width = 1,                    .awvalid
		.s0_axi4lite_awready (axil_driver_0_axil_driver_axi4_lite_awready),           //  output,    width = 1,                    .awready
		.s0_axi4lite_araddr  (axil_driver_0_axil_driver_axi4_lite_araddr),            //   input,   width = 27,                    .araddr
		.s0_axi4lite_arprot  (axil_driver_0_axil_driver_axi4_lite_arprot),            //   input,    width = 3,                    .arprot
		.s0_axi4lite_arvalid (axil_driver_0_axil_driver_axi4_lite_arvalid),           //   input,    width = 1,                    .arvalid
		.s0_axi4lite_arready (axil_driver_0_axil_driver_axi4_lite_arready),           //  output,    width = 1,                    .arready
		.s0_axi4lite_wdata   (axil_driver_0_axil_driver_axi4_lite_wdata),             //   input,   width = 32,                    .wdata
		.s0_axi4lite_wstrb   (axil_driver_0_axil_driver_axi4_lite_wstrb),             //   input,    width = 4,                    .wstrb
		.s0_axi4lite_wvalid  (axil_driver_0_axil_driver_axi4_lite_wvalid),            //   input,    width = 1,                    .wvalid
		.s0_axi4lite_wready  (axil_driver_0_axil_driver_axi4_lite_wready),            //  output,    width = 1,                    .wready
		.s0_axi4lite_bready  (axil_driver_0_axil_driver_axi4_lite_bready),            //   input,    width = 1,                    .bready
		.s0_axi4lite_bresp   (axil_driver_0_axil_driver_axi4_lite_bresp),             //  output,    width = 2,                    .bresp
		.s0_axi4lite_bvalid  (axil_driver_0_axil_driver_axi4_lite_bvalid),            //  output,    width = 1,                    .bvalid
		.s0_axi4lite_rready  (axil_driver_0_axil_driver_axi4_lite_rready),            //   input,    width = 1,                    .rready
		.s0_axi4lite_rdata   (axil_driver_0_axil_driver_axi4_lite_rdata),             //  output,   width = 32,                    .rdata
		.s0_axi4lite_rresp   (axil_driver_0_axil_driver_axi4_lite_rresp),             //  output,    width = 2,                    .rresp
		.s0_axi4lite_rvalid  (axil_driver_0_axil_driver_axi4_lite_rvalid),            //  output,    width = 1,                    .rvalid
		.mem_0_cs            (emif_io96b_lpddr4_0_mem_0_mem_cs),                      //  output,    width = 1,               mem_0.mem_cs
		.mem_0_ca            (emif_io96b_lpddr4_0_mem_0_mem_ca),                      //  output,    width = 6,                    .mem_ca
		.mem_0_cke           (emif_io96b_lpddr4_0_mem_0_mem_cke),                     //  output,    width = 1,                    .mem_cke
		.mem_0_dq            (emif_io96b_lpddr4_0_mem_0_mem_dq),                      //   inout,   width = 32,                    .mem_dq
		.mem_0_dqs_t         (emif_io96b_lpddr4_0_mem_0_mem_dqs_t),                   //   inout,    width = 4,                    .mem_dqs_t
		.mem_0_dqs_c         (emif_io96b_lpddr4_0_mem_0_mem_dqs_c),                   //   inout,    width = 4,                    .mem_dqs_c
		.mem_0_dmi           (emif_io96b_lpddr4_0_mem_0_mem_dmi),                     //   inout,    width = 4,                    .mem_dmi
		.mem_0_ck_t          (emif_io96b_lpddr4_0_mem_ck_0_mem_ck_t),                 //  output,    width = 1,            mem_ck_0.mem_ck_t
		.mem_0_ck_c          (emif_io96b_lpddr4_0_mem_ck_0_mem_ck_c),                 //  output,    width = 1,                    .mem_ck_c
		.mem_0_reset_n       (emif_io96b_lpddr4_0_mem_reset_n_mem_reset_n),           //  output,    width = 1,         mem_reset_n.mem_reset_n
		.oct_rzqin_0         (mem_oct_0_oct_rzqin),                                   //   input,    width = 1,               oct_0.oct_rzqin
		.ref_clk             (ref_clk_source_0_clk_clk)                               //   input,    width = 1,             ref_clk.clk
	);

	ed_sim_mem mem (
		.mem_cke_0     (emif_io96b_lpddr4_0_mem_0_mem_cke),           //   input,   width = 1,       mem_0.mem_cke
		.mem_cs_0      (emif_io96b_lpddr4_0_mem_0_mem_cs),            //   input,   width = 1,            .mem_cs
		.mem_ca_0      (emif_io96b_lpddr4_0_mem_0_mem_ca),            //   input,   width = 6,            .mem_ca
		.mem_dq_0      (emif_io96b_lpddr4_0_mem_0_mem_dq),            //   inout,  width = 32,            .mem_dq
		.mem_dqs_t_0   (emif_io96b_lpddr4_0_mem_0_mem_dqs_t),         //   inout,   width = 4,            .mem_dqs_t
		.mem_dqs_c_0   (emif_io96b_lpddr4_0_mem_0_mem_dqs_c),         //   inout,   width = 4,            .mem_dqs_c
		.mem_dmi_0     (emif_io96b_lpddr4_0_mem_0_mem_dmi),           //   inout,   width = 4,            .mem_dmi
		.mem_ck_t_0    (emif_io96b_lpddr4_0_mem_ck_0_mem_ck_t),       //   input,   width = 1,    mem_ck_0.mem_ck_t
		.mem_ck_c_0    (emif_io96b_lpddr4_0_mem_ck_0_mem_ck_c),       //   input,   width = 1,            .mem_ck_c
		.oct_rzqin_0   (mem_oct_0_oct_rzqin),                         //  output,   width = 1,       oct_0.oct_rzqin
		.mem_reset_n_0 (emif_io96b_lpddr4_0_mem_reset_n_mem_reset_n)  //   input,   width = 1, mem_reset_n.mem_reset_n
	);

	ed_sim_ref_clk_source_0 ref_clk_source_0 (
		.clk (ref_clk_source_0_clk_clk)  //  output,  width = 1, clk.clk
	);

	ed_sim_reset_handler reset_handler (
		.reset_n_0   (~rrip_ninit_done_reset),          //   input,  width = 1,   reset_n_0.reset_n
		.conduit_0   (user_pll_locked_export),          //   input,  width = 1,   conduit_0.export
		.clk         (user_pll_outclk0_clk),            //   input,  width = 1,         clk.clk
		.reset_out_n (reset_handler_reset_n_out_reset)  //  output,  width = 1, reset_n_out.reset_n
	);

	ed_sim_rrip rrip (
		.ninit_done (rrip_ninit_done_reset)  //  output,  width = 1, ninit_done.reset
	);

	ed_sim_traffic_generator traffic_generator (
		.remote_intf_clk              (user_pll_outclk1_clk),                   //   input,    width = 1,   remote_intf_clk.clk
		.remote_intf_reset_n          (reset_handler_reset_n_out_reset),        //   input,    width = 1, remote_intf_reset.reset_n
		.master_jtag_reset_jtag_reset (),                                       //  output,    width = 1,        jtag_reset.reset
		.driver0_axi4_awready         (traffic_generator_driver0_axi4_awready), //   input,    width = 1,      driver0_axi4.awready
		.driver0_axi4_awvalid         (traffic_generator_driver0_axi4_awvalid), //  output,    width = 1,                  .awvalid
		.driver0_axi4_awid            (traffic_generator_driver0_axi4_awid),    //  output,    width = 7,                  .awid
		.driver0_axi4_awaddr          (traffic_generator_driver0_axi4_awaddr),  //  output,   width = 32,                  .awaddr
		.driver0_axi4_awlen           (traffic_generator_driver0_axi4_awlen),   //  output,    width = 8,                  .awlen
		.driver0_axi4_awsize          (traffic_generator_driver0_axi4_awsize),  //  output,    width = 3,                  .awsize
		.driver0_axi4_awburst         (traffic_generator_driver0_axi4_awburst), //  output,    width = 2,                  .awburst
		.driver0_axi4_awlock          (traffic_generator_driver0_axi4_awlock),  //  output,    width = 1,                  .awlock
		.driver0_axi4_awcache         (traffic_generator_driver0_axi4_awcache), //  output,    width = 4,                  .awcache
		.driver0_axi4_awprot          (traffic_generator_driver0_axi4_awprot),  //  output,    width = 3,                  .awprot
		.driver0_axi4_awuser          (traffic_generator_driver0_axi4_awuser),  //  output,    width = 1,                  .awuser
		.driver0_axi4_arready         (traffic_generator_driver0_axi4_arready), //   input,    width = 1,                  .arready
		.driver0_axi4_arvalid         (traffic_generator_driver0_axi4_arvalid), //  output,    width = 1,                  .arvalid
		.driver0_axi4_arid            (traffic_generator_driver0_axi4_arid),    //  output,    width = 7,                  .arid
		.driver0_axi4_araddr          (traffic_generator_driver0_axi4_araddr),  //  output,   width = 32,                  .araddr
		.driver0_axi4_arlen           (traffic_generator_driver0_axi4_arlen),   //  output,    width = 8,                  .arlen
		.driver0_axi4_arsize          (traffic_generator_driver0_axi4_arsize),  //  output,    width = 3,                  .arsize
		.driver0_axi4_arburst         (traffic_generator_driver0_axi4_arburst), //  output,    width = 2,                  .arburst
		.driver0_axi4_arlock          (traffic_generator_driver0_axi4_arlock),  //  output,    width = 1,                  .arlock
		.driver0_axi4_arcache         (traffic_generator_driver0_axi4_arcache), //  output,    width = 4,                  .arcache
		.driver0_axi4_arprot          (traffic_generator_driver0_axi4_arprot),  //  output,    width = 3,                  .arprot
		.driver0_axi4_aruser          (traffic_generator_driver0_axi4_aruser),  //  output,    width = 1,                  .aruser
		.driver0_axi4_wready          (traffic_generator_driver0_axi4_wready),  //   input,    width = 1,                  .wready
		.driver0_axi4_wvalid          (traffic_generator_driver0_axi4_wvalid),  //  output,    width = 1,                  .wvalid
		.driver0_axi4_wdata           (traffic_generator_driver0_axi4_wdata),   //  output,  width = 256,                  .wdata
		.driver0_axi4_wstrb           (traffic_generator_driver0_axi4_wstrb),   //  output,   width = 32,                  .wstrb
		.driver0_axi4_wlast           (traffic_generator_driver0_axi4_wlast),   //  output,    width = 1,                  .wlast
		.driver0_axi4_bready          (traffic_generator_driver0_axi4_bready),  //  output,    width = 1,                  .bready
		.driver0_axi4_bvalid          (traffic_generator_driver0_axi4_bvalid),  //   input,    width = 1,                  .bvalid
		.driver0_axi4_bid             (traffic_generator_driver0_axi4_bid),     //   input,    width = 7,                  .bid
		.driver0_axi4_bresp           (traffic_generator_driver0_axi4_bresp),   //   input,    width = 2,                  .bresp
		.driver0_axi4_rready          (traffic_generator_driver0_axi4_rready),  //  output,    width = 1,                  .rready
		.driver0_axi4_rvalid          (traffic_generator_driver0_axi4_rvalid),  //   input,    width = 1,                  .rvalid
		.driver0_axi4_rid             (traffic_generator_driver0_axi4_rid),     //   input,    width = 7,                  .rid
		.driver0_axi4_rdata           (traffic_generator_driver0_axi4_rdata),   //   input,  width = 256,                  .rdata
		.driver0_axi4_rresp           (traffic_generator_driver0_axi4_rresp),   //   input,    width = 2,                  .rresp
		.driver0_axi4_rlast           (traffic_generator_driver0_axi4_rlast),   //   input,    width = 1,                  .rlast
		.driver0_clk                  (user_pll_outclk0_clk),                   //   input,    width = 1,       driver0_clk.clk
		.driver0_reset_n              (axil_driver_0_cal_done_rst_n_reset)      //   input,    width = 1,     driver0_reset.reset_n
	);

	ed_sim_user_pll user_pll (
		.refclk   (async_clk_source_clk_clk), //   input,  width = 1,  refclk.clk
		.locked   (user_pll_locked_export),   //  output,  width = 1,  locked.export
		.rst      (rrip_ninit_done_reset),    //   input,  width = 1,   reset.reset
		.outclk_0 (user_pll_outclk0_clk),     //  output,  width = 1, outclk0.clk
		.outclk_1 (user_pll_outclk1_clk)      //  output,  width = 1, outclk1.clk
	);

	ed_sim_altera_mm_interconnect_1920_h43vqey mm_interconnect_1 (
		.traffic_generator_driver0_axi4_awid                                             (traffic_generator_driver0_axi4_awid),                   //   input,    width = 7,                                            traffic_generator_driver0_axi4.awid
		.traffic_generator_driver0_axi4_awaddr                                           (traffic_generator_driver0_axi4_awaddr),                 //   input,   width = 32,                                                                          .awaddr
		.traffic_generator_driver0_axi4_awlen                                            (traffic_generator_driver0_axi4_awlen),                  //   input,    width = 8,                                                                          .awlen
		.traffic_generator_driver0_axi4_awsize                                           (traffic_generator_driver0_axi4_awsize),                 //   input,    width = 3,                                                                          .awsize
		.traffic_generator_driver0_axi4_awburst                                          (traffic_generator_driver0_axi4_awburst),                //   input,    width = 2,                                                                          .awburst
		.traffic_generator_driver0_axi4_awlock                                           (traffic_generator_driver0_axi4_awlock),                 //   input,    width = 1,                                                                          .awlock
		.traffic_generator_driver0_axi4_awcache                                          (traffic_generator_driver0_axi4_awcache),                //   input,    width = 4,                                                                          .awcache
		.traffic_generator_driver0_axi4_awprot                                           (traffic_generator_driver0_axi4_awprot),                 //   input,    width = 3,                                                                          .awprot
		.traffic_generator_driver0_axi4_awuser                                           (traffic_generator_driver0_axi4_awuser),                 //   input,    width = 1,                                                                          .awuser
		.traffic_generator_driver0_axi4_awvalid                                          (traffic_generator_driver0_axi4_awvalid),                //   input,    width = 1,                                                                          .awvalid
		.traffic_generator_driver0_axi4_awready                                          (traffic_generator_driver0_axi4_awready),                //  output,    width = 1,                                                                          .awready
		.traffic_generator_driver0_axi4_wdata                                            (traffic_generator_driver0_axi4_wdata),                  //   input,  width = 256,                                                                          .wdata
		.traffic_generator_driver0_axi4_wstrb                                            (traffic_generator_driver0_axi4_wstrb),                  //   input,   width = 32,                                                                          .wstrb
		.traffic_generator_driver0_axi4_wlast                                            (traffic_generator_driver0_axi4_wlast),                  //   input,    width = 1,                                                                          .wlast
		.traffic_generator_driver0_axi4_wvalid                                           (traffic_generator_driver0_axi4_wvalid),                 //   input,    width = 1,                                                                          .wvalid
		.traffic_generator_driver0_axi4_wready                                           (traffic_generator_driver0_axi4_wready),                 //  output,    width = 1,                                                                          .wready
		.traffic_generator_driver0_axi4_bid                                              (traffic_generator_driver0_axi4_bid),                    //  output,    width = 7,                                                                          .bid
		.traffic_generator_driver0_axi4_bresp                                            (traffic_generator_driver0_axi4_bresp),                  //  output,    width = 2,                                                                          .bresp
		.traffic_generator_driver0_axi4_bvalid                                           (traffic_generator_driver0_axi4_bvalid),                 //  output,    width = 1,                                                                          .bvalid
		.traffic_generator_driver0_axi4_bready                                           (traffic_generator_driver0_axi4_bready),                 //   input,    width = 1,                                                                          .bready
		.traffic_generator_driver0_axi4_arid                                             (traffic_generator_driver0_axi4_arid),                   //   input,    width = 7,                                                                          .arid
		.traffic_generator_driver0_axi4_araddr                                           (traffic_generator_driver0_axi4_araddr),                 //   input,   width = 32,                                                                          .araddr
		.traffic_generator_driver0_axi4_arlen                                            (traffic_generator_driver0_axi4_arlen),                  //   input,    width = 8,                                                                          .arlen
		.traffic_generator_driver0_axi4_arsize                                           (traffic_generator_driver0_axi4_arsize),                 //   input,    width = 3,                                                                          .arsize
		.traffic_generator_driver0_axi4_arburst                                          (traffic_generator_driver0_axi4_arburst),                //   input,    width = 2,                                                                          .arburst
		.traffic_generator_driver0_axi4_arlock                                           (traffic_generator_driver0_axi4_arlock),                 //   input,    width = 1,                                                                          .arlock
		.traffic_generator_driver0_axi4_arcache                                          (traffic_generator_driver0_axi4_arcache),                //   input,    width = 4,                                                                          .arcache
		.traffic_generator_driver0_axi4_arprot                                           (traffic_generator_driver0_axi4_arprot),                 //   input,    width = 3,                                                                          .arprot
		.traffic_generator_driver0_axi4_aruser                                           (traffic_generator_driver0_axi4_aruser),                 //   input,    width = 1,                                                                          .aruser
		.traffic_generator_driver0_axi4_arvalid                                          (traffic_generator_driver0_axi4_arvalid),                //   input,    width = 1,                                                                          .arvalid
		.traffic_generator_driver0_axi4_arready                                          (traffic_generator_driver0_axi4_arready),                //  output,    width = 1,                                                                          .arready
		.traffic_generator_driver0_axi4_rid                                              (traffic_generator_driver0_axi4_rid),                    //  output,    width = 7,                                                                          .rid
		.traffic_generator_driver0_axi4_rdata                                            (traffic_generator_driver0_axi4_rdata),                  //  output,  width = 256,                                                                          .rdata
		.traffic_generator_driver0_axi4_rresp                                            (traffic_generator_driver0_axi4_rresp),                  //  output,    width = 2,                                                                          .rresp
		.traffic_generator_driver0_axi4_rlast                                            (traffic_generator_driver0_axi4_rlast),                  //  output,    width = 1,                                                                          .rlast
		.traffic_generator_driver0_axi4_rvalid                                           (traffic_generator_driver0_axi4_rvalid),                 //  output,    width = 1,                                                                          .rvalid
		.traffic_generator_driver0_axi4_rready                                           (traffic_generator_driver0_axi4_rready),                 //   input,    width = 1,                                                                          .rready
		.emif_io96b_lpddr4_0_s0_axi4_awid                                                (mm_interconnect_1_emif_io96b_lpddr4_0_s0_axi4_awid),    //  output,    width = 7,                                               emif_io96b_lpddr4_0_s0_axi4.awid
		.emif_io96b_lpddr4_0_s0_axi4_awaddr                                              (mm_interconnect_1_emif_io96b_lpddr4_0_s0_axi4_awaddr),  //  output,   width = 32,                                                                          .awaddr
		.emif_io96b_lpddr4_0_s0_axi4_awlen                                               (mm_interconnect_1_emif_io96b_lpddr4_0_s0_axi4_awlen),   //  output,    width = 8,                                                                          .awlen
		.emif_io96b_lpddr4_0_s0_axi4_awsize                                              (mm_interconnect_1_emif_io96b_lpddr4_0_s0_axi4_awsize),  //  output,    width = 3,                                                                          .awsize
		.emif_io96b_lpddr4_0_s0_axi4_awburst                                             (mm_interconnect_1_emif_io96b_lpddr4_0_s0_axi4_awburst), //  output,    width = 2,                                                                          .awburst
		.emif_io96b_lpddr4_0_s0_axi4_awlock                                              (mm_interconnect_1_emif_io96b_lpddr4_0_s0_axi4_awlock),  //  output,    width = 1,                                                                          .awlock
		.emif_io96b_lpddr4_0_s0_axi4_awprot                                              (mm_interconnect_1_emif_io96b_lpddr4_0_s0_axi4_awprot),  //  output,    width = 3,                                                                          .awprot
		.emif_io96b_lpddr4_0_s0_axi4_awuser                                              (mm_interconnect_1_emif_io96b_lpddr4_0_s0_axi4_awuser),  //  output,   width = 14,                                                                          .awuser
		.emif_io96b_lpddr4_0_s0_axi4_awqos                                               (mm_interconnect_1_emif_io96b_lpddr4_0_s0_axi4_awqos),   //  output,    width = 4,                                                                          .awqos
		.emif_io96b_lpddr4_0_s0_axi4_awvalid                                             (mm_interconnect_1_emif_io96b_lpddr4_0_s0_axi4_awvalid), //  output,    width = 1,                                                                          .awvalid
		.emif_io96b_lpddr4_0_s0_axi4_awready                                             (mm_interconnect_1_emif_io96b_lpddr4_0_s0_axi4_awready), //   input,    width = 1,                                                                          .awready
		.emif_io96b_lpddr4_0_s0_axi4_wdata                                               (mm_interconnect_1_emif_io96b_lpddr4_0_s0_axi4_wdata),   //  output,  width = 256,                                                                          .wdata
		.emif_io96b_lpddr4_0_s0_axi4_wstrb                                               (mm_interconnect_1_emif_io96b_lpddr4_0_s0_axi4_wstrb),   //  output,   width = 32,                                                                          .wstrb
		.emif_io96b_lpddr4_0_s0_axi4_wlast                                               (mm_interconnect_1_emif_io96b_lpddr4_0_s0_axi4_wlast),   //  output,    width = 1,                                                                          .wlast
		.emif_io96b_lpddr4_0_s0_axi4_wvalid                                              (mm_interconnect_1_emif_io96b_lpddr4_0_s0_axi4_wvalid),  //  output,    width = 1,                                                                          .wvalid
		.emif_io96b_lpddr4_0_s0_axi4_wuser                                               (mm_interconnect_1_emif_io96b_lpddr4_0_s0_axi4_wuser),   //  output,   width = 32,                                                                          .wuser
		.emif_io96b_lpddr4_0_s0_axi4_wready                                              (mm_interconnect_1_emif_io96b_lpddr4_0_s0_axi4_wready),  //   input,    width = 1,                                                                          .wready
		.emif_io96b_lpddr4_0_s0_axi4_bid                                                 (mm_interconnect_1_emif_io96b_lpddr4_0_s0_axi4_bid),     //   input,    width = 7,                                                                          .bid
		.emif_io96b_lpddr4_0_s0_axi4_bresp                                               (mm_interconnect_1_emif_io96b_lpddr4_0_s0_axi4_bresp),   //   input,    width = 2,                                                                          .bresp
		.emif_io96b_lpddr4_0_s0_axi4_bvalid                                              (mm_interconnect_1_emif_io96b_lpddr4_0_s0_axi4_bvalid),  //   input,    width = 1,                                                                          .bvalid
		.emif_io96b_lpddr4_0_s0_axi4_bready                                              (mm_interconnect_1_emif_io96b_lpddr4_0_s0_axi4_bready),  //  output,    width = 1,                                                                          .bready
		.emif_io96b_lpddr4_0_s0_axi4_arid                                                (mm_interconnect_1_emif_io96b_lpddr4_0_s0_axi4_arid),    //  output,    width = 7,                                                                          .arid
		.emif_io96b_lpddr4_0_s0_axi4_araddr                                              (mm_interconnect_1_emif_io96b_lpddr4_0_s0_axi4_araddr),  //  output,   width = 32,                                                                          .araddr
		.emif_io96b_lpddr4_0_s0_axi4_arlen                                               (mm_interconnect_1_emif_io96b_lpddr4_0_s0_axi4_arlen),   //  output,    width = 8,                                                                          .arlen
		.emif_io96b_lpddr4_0_s0_axi4_arsize                                              (mm_interconnect_1_emif_io96b_lpddr4_0_s0_axi4_arsize),  //  output,    width = 3,                                                                          .arsize
		.emif_io96b_lpddr4_0_s0_axi4_arburst                                             (mm_interconnect_1_emif_io96b_lpddr4_0_s0_axi4_arburst), //  output,    width = 2,                                                                          .arburst
		.emif_io96b_lpddr4_0_s0_axi4_arlock                                              (mm_interconnect_1_emif_io96b_lpddr4_0_s0_axi4_arlock),  //  output,    width = 1,                                                                          .arlock
		.emif_io96b_lpddr4_0_s0_axi4_arprot                                              (mm_interconnect_1_emif_io96b_lpddr4_0_s0_axi4_arprot),  //  output,    width = 3,                                                                          .arprot
		.emif_io96b_lpddr4_0_s0_axi4_aruser                                              (mm_interconnect_1_emif_io96b_lpddr4_0_s0_axi4_aruser),  //  output,   width = 14,                                                                          .aruser
		.emif_io96b_lpddr4_0_s0_axi4_arqos                                               (mm_interconnect_1_emif_io96b_lpddr4_0_s0_axi4_arqos),   //  output,    width = 4,                                                                          .arqos
		.emif_io96b_lpddr4_0_s0_axi4_arvalid                                             (mm_interconnect_1_emif_io96b_lpddr4_0_s0_axi4_arvalid), //  output,    width = 1,                                                                          .arvalid
		.emif_io96b_lpddr4_0_s0_axi4_arready                                             (mm_interconnect_1_emif_io96b_lpddr4_0_s0_axi4_arready), //   input,    width = 1,                                                                          .arready
		.emif_io96b_lpddr4_0_s0_axi4_rid                                                 (mm_interconnect_1_emif_io96b_lpddr4_0_s0_axi4_rid),     //   input,    width = 7,                                                                          .rid
		.emif_io96b_lpddr4_0_s0_axi4_rdata                                               (mm_interconnect_1_emif_io96b_lpddr4_0_s0_axi4_rdata),   //   input,  width = 256,                                                                          .rdata
		.emif_io96b_lpddr4_0_s0_axi4_rresp                                               (mm_interconnect_1_emif_io96b_lpddr4_0_s0_axi4_rresp),   //   input,    width = 2,                                                                          .rresp
		.emif_io96b_lpddr4_0_s0_axi4_rlast                                               (mm_interconnect_1_emif_io96b_lpddr4_0_s0_axi4_rlast),   //   input,    width = 1,                                                                          .rlast
		.emif_io96b_lpddr4_0_s0_axi4_rvalid                                              (mm_interconnect_1_emif_io96b_lpddr4_0_s0_axi4_rvalid),  //   input,    width = 1,                                                                          .rvalid
		.emif_io96b_lpddr4_0_s0_axi4_rready                                              (mm_interconnect_1_emif_io96b_lpddr4_0_s0_axi4_rready),  //  output,    width = 1,                                                                          .rready
		.emif_io96b_lpddr4_0_s0_axi4_ruser                                               (mm_interconnect_1_emif_io96b_lpddr4_0_s0_axi4_ruser),   //   input,   width = 32,                                                                          .ruser
		.traffic_generator_driver0_axi4_translator_clk_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                    //   input,    width = 1, traffic_generator_driver0_axi4_translator_clk_reset_reset_bridge_in_reset.reset
		.emif_io96b_lpddr4_0_s0_axi4_translator_clk_reset_reset_bridge_in_reset_reset    (rst_controller_002_reset_out_reset),                    //   input,    width = 1,    emif_io96b_lpddr4_0_s0_axi4_translator_clk_reset_reset_bridge_in_reset.reset
		.user_pll_outclk0_clk                                                            (user_pll_outclk0_clk)                                   //   input,    width = 1,                                                          user_pll_outclk0.clk
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_handler_reset_n_out_reset), //   input,  width = 1, reset_in0.reset
		.clk            (user_pll_outclk1_clk),             //   input,  width = 1,       clk.clk
		.reset_out      (rst_controller_reset_out_reset),   //  output,  width = 1, reset_out.reset
		.reset_req      (),                                 // (terminated),                       
		.reset_req_in0  (1'b0),                             // (terminated),                       
		.reset_in1      (1'b0),                             // (terminated),                       
		.reset_req_in1  (1'b0),                             // (terminated),                       
		.reset_in2      (1'b0),                             // (terminated),                       
		.reset_req_in2  (1'b0),                             // (terminated),                       
		.reset_in3      (1'b0),                             // (terminated),                       
		.reset_req_in3  (1'b0),                             // (terminated),                       
		.reset_in4      (1'b0),                             // (terminated),                       
		.reset_req_in4  (1'b0),                             // (terminated),                       
		.reset_in5      (1'b0),                             // (terminated),                       
		.reset_req_in5  (1'b0),                             // (terminated),                       
		.reset_in6      (1'b0),                             // (terminated),                       
		.reset_req_in6  (1'b0),                             // (terminated),                       
		.reset_in7      (1'b0),                             // (terminated),                       
		.reset_req_in7  (1'b0),                             // (terminated),                       
		.reset_in8      (1'b0),                             // (terminated),                       
		.reset_req_in8  (1'b0),                             // (terminated),                       
		.reset_in9      (1'b0),                             // (terminated),                       
		.reset_req_in9  (1'b0),                             // (terminated),                       
		.reset_in10     (1'b0),                             // (terminated),                       
		.reset_req_in10 (1'b0),                             // (terminated),                       
		.reset_in11     (1'b0),                             // (terminated),                       
		.reset_req_in11 (1'b0),                             // (terminated),                       
		.reset_in12     (1'b0),                             // (terminated),                       
		.reset_req_in12 (1'b0),                             // (terminated),                       
		.reset_in13     (1'b0),                             // (terminated),                       
		.reset_req_in13 (1'b0),                             // (terminated),                       
		.reset_in14     (1'b0),                             // (terminated),                       
		.reset_req_in14 (1'b0),                             // (terminated),                       
		.reset_in15     (1'b0),                             // (terminated),                       
		.reset_req_in15 (1'b0)                              // (terminated),                       
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("both"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~axil_driver_0_cal_done_rst_n_reset), //   input,  width = 1, reset_in0.reset
		.clk            (user_pll_outclk0_clk),                //   input,  width = 1,       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),  //  output,  width = 1, reset_out.reset
		.reset_req      (),                                    // (terminated),                       
		.reset_req_in0  (1'b0),                                // (terminated),                       
		.reset_in1      (1'b0),                                // (terminated),                       
		.reset_req_in1  (1'b0),                                // (terminated),                       
		.reset_in2      (1'b0),                                // (terminated),                       
		.reset_req_in2  (1'b0),                                // (terminated),                       
		.reset_in3      (1'b0),                                // (terminated),                       
		.reset_req_in3  (1'b0),                                // (terminated),                       
		.reset_in4      (1'b0),                                // (terminated),                       
		.reset_req_in4  (1'b0),                                // (terminated),                       
		.reset_in5      (1'b0),                                // (terminated),                       
		.reset_req_in5  (1'b0),                                // (terminated),                       
		.reset_in6      (1'b0),                                // (terminated),                       
		.reset_req_in6  (1'b0),                                // (terminated),                       
		.reset_in7      (1'b0),                                // (terminated),                       
		.reset_req_in7  (1'b0),                                // (terminated),                       
		.reset_in8      (1'b0),                                // (terminated),                       
		.reset_req_in8  (1'b0),                                // (terminated),                       
		.reset_in9      (1'b0),                                // (terminated),                       
		.reset_req_in9  (1'b0),                                // (terminated),                       
		.reset_in10     (1'b0),                                // (terminated),                       
		.reset_req_in10 (1'b0),                                // (terminated),                       
		.reset_in11     (1'b0),                                // (terminated),                       
		.reset_req_in11 (1'b0),                                // (terminated),                       
		.reset_in12     (1'b0),                                // (terminated),                       
		.reset_req_in12 (1'b0),                                // (terminated),                       
		.reset_in13     (1'b0),                                // (terminated),                       
		.reset_req_in13 (1'b0),                                // (terminated),                       
		.reset_in14     (1'b0),                                // (terminated),                       
		.reset_req_in14 (1'b0),                                // (terminated),                       
		.reset_in15     (1'b0),                                // (terminated),                       
		.reset_req_in15 (1'b0)                                 // (terminated),                       
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("both"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~emif_io96b_lpddr4_0_s0_axi4_ctrl_ready_reset), //   input,  width = 1, reset_in0.reset
		.clk            (user_pll_outclk0_clk),                          //   input,  width = 1,       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset),            //  output,  width = 1, reset_out.reset
		.reset_req      (),                                              // (terminated),                       
		.reset_req_in0  (1'b0),                                          // (terminated),                       
		.reset_in1      (1'b0),                                          // (terminated),                       
		.reset_req_in1  (1'b0),                                          // (terminated),                       
		.reset_in2      (1'b0),                                          // (terminated),                       
		.reset_req_in2  (1'b0),                                          // (terminated),                       
		.reset_in3      (1'b0),                                          // (terminated),                       
		.reset_req_in3  (1'b0),                                          // (terminated),                       
		.reset_in4      (1'b0),                                          // (terminated),                       
		.reset_req_in4  (1'b0),                                          // (terminated),                       
		.reset_in5      (1'b0),                                          // (terminated),                       
		.reset_req_in5  (1'b0),                                          // (terminated),                       
		.reset_in6      (1'b0),                                          // (terminated),                       
		.reset_req_in6  (1'b0),                                          // (terminated),                       
		.reset_in7      (1'b0),                                          // (terminated),                       
		.reset_req_in7  (1'b0),                                          // (terminated),                       
		.reset_in8      (1'b0),                                          // (terminated),                       
		.reset_req_in8  (1'b0),                                          // (terminated),                       
		.reset_in9      (1'b0),                                          // (terminated),                       
		.reset_req_in9  (1'b0),                                          // (terminated),                       
		.reset_in10     (1'b0),                                          // (terminated),                       
		.reset_req_in10 (1'b0),                                          // (terminated),                       
		.reset_in11     (1'b0),                                          // (terminated),                       
		.reset_req_in11 (1'b0),                                          // (terminated),                       
		.reset_in12     (1'b0),                                          // (terminated),                       
		.reset_req_in12 (1'b0),                                          // (terminated),                       
		.reset_in13     (1'b0),                                          // (terminated),                       
		.reset_req_in13 (1'b0),                                          // (terminated),                       
		.reset_in14     (1'b0),                                          // (terminated),                       
		.reset_req_in14 (1'b0),                                          // (terminated),                       
		.reset_in15     (1'b0),                                          // (terminated),                       
		.reset_req_in15 (1'b0)                                           // (terminated),                       
	);

endmodule
