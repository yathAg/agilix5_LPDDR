module ed_sim (
	);
endmodule

